library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;
---------------------------------------------------------------------------------------------------------------------------------
-- ENTITY DECLARATION
---------------------------------------------------------------------------------------------------------------------------------
entity frame_vga is
    Port (  -- CLOCK 
            FRM_i_CLK_100M  :   in  std_logic;
            FRM_i_CLK_25M   :   in  std_logic;
            -- IN DELAY
            FRM_i_DONE      :   in  std_logic                    ;
            -- IN GAMELOGIC 
            FRM_i_CURS_X    :   in  std_logic_vector( 3 downto 0);
            FRM_i_CURS_Y    :   in  std_logic_vector( 3 downto 0);
            FRM_i_PIECE     :   in  std_logic_vector( 9 downto 0);
            -- INPUT DA VGA 
            FRM_i_ON_STATE  :   in  std_logic                    ;
            FRM_i_V_CNT     :   in  std_logic_vector(10 downto 0);
            FRM_i_H_CNT     :   in  std_logic_vector(10 downto 0);            
            -- OUT DELAY
            FRM_o_DELAY_MS  :   out std_logic_vector(11 downto 0);
            FRM_o_DELAY_EN  :   out std_logic                    ;
            -- OUTPUT A VGA
            FRM_o_R         :   out std_logic_vector( 3 downto 0);
            FRM_o_G         :   out std_logic_vector( 3 downto 0);
            FRM_o_B         :   out std_logic_vector( 3 downto 0);
            -- OUTPUT A GAME_LOGIC
            FRM_o_ACK       :   out std_logic                    );
end frame_vga;
---------------------------------------------------------------------------------------------------------------------------------
-- ARCHITECTURE DECLARATION                                                                                                            
---------------------------------------------------------------------------------------------------------------------------------
architecture Behavioral of frame_vga is
---------------------------------------------------------------------------------------------------------------------------------
-- TYPE DECLARATION                                                                                                      
--------------------------------------------------------------------------------------------------------------------------------- 
    type tp_cella is array(0 to 19, 0 to 19) of std_logic_vector(11 downto 0);
    type tp_stato is (  IDLE    ,
                        LAMP_ON ,
                        LAMP_OFF,
                        WAIT1   ,
                        WAIT2   ,
                        WAIT3   );
---------------------------------------------------------------------------------------------------------------------------------
-- CONSTANT DECLARATION                                                                                                       
---------------------------------------------------------------------------------------------------------------------------------
    -- Bianco
    constant empty_L : tp_cella := ((x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF"),
                                    (x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF"),
                                    (x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF"),
                                    (x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF"),
                                    (x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF"),
                                    (x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF"),
                                    (x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF"),
                                    (x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF"),
                                    (x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF"),
                                    (x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF"),
                                    (x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF"),
                                    (x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF"),
                                    (x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF"),
                                    (x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF"),
                                    (x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF"),
                                    (x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF"),
                                    (x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF"),
                                    (x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF"),
                                    (x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF"),
                                    (x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF", x"FFF"));
    constant pawn_L : tp_cella :=  ((x"F00", x"F00", x"F00", x"F00", x"F00", x"F00", x"F00", x"F00", x"F00", x"F00", x"F00", x"F00", x"F00", x"F00", x"F00", x"F00", x"F00", x"F00", x"F00", x"F00"),
                                    (x"F00", x"444", x"444", x"444", x"444", x"444", x"444", x"444", x"F00", x"F00", x"F00", x"444", x"444", x"444", x"444", x"444", x"444", x"444", x"F00", x"F00"),
                                    (x"F00", x"444", x"444", x"444", x"444", x"444", x"444", x"444", x"F00", x"F00", x"F00", x"444", x"444", x"444", x"444", x"444", x"444", x"444", x"F00", x"F00"),
                                    (x"F00", x"444", x"444", x"444", x"444", x"444", x"444", x"444", x"F00", x"F00", x"F00", x"444", x"444", x"444", x"444", x"444", x"444", x"444", x"F00", x"F00"),
                                    (x"F00", x"444", x"444", x"444", x"444", x"444", x"444", x"444", x"F00", x"F00", x"F00", x"444", x"444", x"444", x"444", x"444", x"444", x"444", x"F00", x"F00"),
                                    (x"F00", x"444", x"444", x"444", x"444", x"444", x"444", x"444", x"F00", x"F00", x"F00", x"444", x"444", x"444", x"444", x"444", x"444", x"444", x"F00", x"F00"),
                                    (x"F00", x"444", x"444", x"444", x"444", x"444", x"444", x"444", x"F00", x"F00", x"F00", x"444", x"444", x"444", x"444", x"444", x"444", x"444", x"F00", x"F00"),
                                    (x"F00", x"444", x"444", x"444", x"444", x"444", x"444", x"444", x"F00", x"F00", x"F00", x"444", x"444", x"444", x"444", x"444", x"444", x"444", x"F00", x"F00"),
                                    (x"F00", x"444", x"444", x"444", x"444", x"444", x"444", x"444", x"F00", x"F00", x"F00", x"444", x"444", x"444", x"444", x"444", x"444", x"444", x"F00", x"F00"),
                                    (x"F00", x"444", x"444", x"444", x"444", x"444", x"444", x"444", x"F00", x"F00", x"F00", x"444", x"444", x"444", x"444", x"444", x"444", x"444", x"F00", x"F00"),
                                    (x"F00", x"444", x"444", x"444", x"444", x"444", x"444", x"444", x"F00", x"F00", x"F00", x"444", x"444", x"444", x"444", x"444", x"444", x"444", x"F00", x"F00"),
                                    (x"F00", x"444", x"444", x"444", x"444", x"444", x"444", x"444", x"F00", x"F00", x"F00", x"444", x"444", x"444", x"444", x"444", x"444", x"444", x"F00", x"F00"),
                                    (x"F00", x"444", x"444", x"444", x"444", x"444", x"444", x"444", x"F00", x"F00", x"F00", x"444", x"444", x"444", x"444", x"444", x"444", x"444", x"F00", x"F00"),
                                    (x"F00", x"444", x"444", x"444", x"444", x"444", x"444", x"444", x"F00", x"F00", x"F00", x"444", x"444", x"444", x"444", x"444", x"444", x"444", x"F00", x"F00"),
                                    (x"F00", x"444", x"444", x"444", x"444", x"444", x"444", x"F00", x"F00", x"F00", x"F00", x"F00", x"444", x"444", x"444", x"444", x"444", x"444", x"F00", x"F00"),
                                    (x"F00", x"444", x"444", x"444", x"444", x"444", x"444", x"F00", x"F00", x"F00", x"F00", x"F00", x"444", x"444", x"444", x"444", x"444", x"444", x"F00", x"F00"),
                                    (x"F00", x"444", x"444", x"444", x"444", x"F00", x"F00", x"F00", x"F00", x"F00", x"F00", x"F00", x"F00", x"F00", x"444", x"444", x"444", x"444", x"F00", x"F00"),
                                    (x"F00", x"444", x"444", x"444", x"F00", x"F00", x"F00", x"F00", x"F00", x"F00", x"F00", x"F00", x"F00", x"F00", x"F00", x"444", x"444", x"444", x"F00", x"F00"),
                                    (x"F00", x"444", x"444", x"F00", x"F00", x"F00", x"F00", x"F00", x"F00", x"F00", x"F00", x"F00", x"F00", x"F00", x"F00", x"F00", x"444", x"444", x"F00", x"F00"),
                                    (x"F00", x"F00", x"F00", x"F00", x"F00", x"F00", x"F00", x"F00", x"F00", x"F00", x"F00", x"F00", x"F00", x"F00", x"F00", x"F00", x"F00", x"F00", x"F00", x"F00"));
    constant king_L : tp_cella :=  ((x"F00", x"F00", x"F00", x"F00", x"F00", x"F00", x"F00", x"F00", x"F00", x"F00", x"F00", x"F00", x"F00", x"F00", x"F00", x"F00", x"F00", x"F00", x"F00", x"F00"),
                                    (x"F00", x"444", x"444", x"444", x"444", x"444", x"444", x"444", x"F00", x"F00", x"444", x"444", x"444", x"444", x"444", x"444", x"444", x"444", x"F00", x"F00"),
                                    (x"F00", x"444", x"444", x"444", x"444", x"444", x"F00", x"F00", x"F00", x"F00", x"F00", x"F00", x"444", x"444", x"444", x"444", x"444", x"444", x"F00", x"F00"),
                                    (x"F00", x"444", x"444", x"444", x"444", x"444", x"F00", x"F00", x"F00", x"F00", x"F00", x"F00", x"444", x"444", x"444", x"444", x"444", x"444", x"F00", x"F00"),
                                    (x"F00", x"444", x"444", x"444", x"444", x"444", x"444", x"444", x"F00", x"F00", x"444", x"444", x"444", x"444", x"444", x"444", x"444", x"444", x"F00", x"F00"),
                                    (x"F00", x"444", x"444", x"444", x"444", x"444", x"444", x"444", x"F00", x"F00", x"444", x"444", x"444", x"444", x"444", x"444", x"444", x"444", x"F00", x"F00"),
                                    (x"F00", x"444", x"444", x"444", x"444", x"444", x"444", x"F00", x"F00", x"F00", x"F00", x"444", x"444", x"444", x"444", x"444", x"444", x"444", x"F00", x"F00"),
                                    (x"F00", x"444", x"444", x"444", x"444", x"444", x"F00", x"F00", x"F00", x"F00", x"F00", x"F00", x"444", x"444", x"444", x"444", x"444", x"444", x"F00", x"F00"),
                                    (x"F00", x"444", x"444", x"444", x"444", x"444", x"F00", x"F00", x"F00", x"F00", x"F00", x"F00", x"444", x"444", x"444", x"444", x"444", x"444", x"F00", x"F00"),
                                    (x"F00", x"444", x"444", x"444", x"444", x"444", x"F00", x"F00", x"F00", x"F00", x"F00", x"F00", x"444", x"444", x"444", x"444", x"444", x"444", x"F00", x"F00"),
                                    (x"F00", x"444", x"444", x"444", x"444", x"F00", x"F00", x"F00", x"F00", x"F00", x"F00", x"F00", x"F00", x"444", x"444", x"444", x"444", x"444", x"F00", x"F00"),
                                    (x"F00", x"444", x"444", x"444", x"444", x"444", x"F00", x"F00", x"F00", x"F00", x"F00", x"F00", x"444", x"444", x"444", x"444", x"444", x"444", x"F00", x"F00"),
                                    (x"F00", x"444", x"444", x"444", x"444", x"444", x"444", x"F00", x"F00", x"F00", x"F00", x"444", x"444", x"444", x"444", x"444", x"444", x"444", x"F00", x"F00"),
                                    (x"F00", x"444", x"444", x"444", x"444", x"444", x"444", x"F00", x"F00", x"F00", x"F00", x"444", x"444", x"444", x"444", x"444", x"444", x"444", x"F00", x"F00"),
                                    (x"F00", x"444", x"444", x"444", x"444", x"444", x"444", x"F00", x"F00", x"F00", x"F00", x"444", x"444", x"444", x"444", x"444", x"444", x"444", x"F00", x"F00"),
                                    (x"F00", x"444", x"444", x"444", x"444", x"444", x"444", x"F00", x"F00", x"F00", x"F00", x"444", x"444", x"444", x"444", x"444", x"444", x"444", x"F00", x"F00"),
                                    (x"F00", x"444", x"444", x"444", x"444", x"444", x"F00", x"F00", x"F00", x"F00", x"F00", x"F00", x"444", x"444", x"444", x"444", x"444", x"444", x"F00", x"F00"),
                                    (x"F00", x"444", x"444", x"444", x"444", x"F00", x"F00", x"F00", x"F00", x"F00", x"F00", x"F00", x"F00", x"444", x"444", x"444", x"444", x"444", x"F00", x"F00"),
                                    (x"F00", x"444", x"444", x"444", x"F00", x"F00", x"F00", x"F00", x"F00", x"F00", x"F00", x"F00", x"F00", x"F00", x"444", x"444", x"444", x"444", x"F00", x"F00"),
                                    (x"F00", x"F00", x"F00", x"F00", x"F00", x"F00", x"F00", x"F00", x"F00", x"F00", x"F00", x"F00", x"F00", x"F00", x"F00", x"F00", x"F00", x"F00", x"F00", x"F00"));
    constant queen_L : tp_cella := ((x"F00", x"F00", x"F00", x"F00", x"F00", x"F00", x"F00", x"F00", x"F00", x"F00", x"F00", x"F00", x"F00", x"F00", x"F00", x"F00", x"F00", x"F00", x"F00", x"F00"),
                                    (x"F00", x"444", x"444", x"444", x"444", x"444", x"444", x"444", x"F00", x"F00", x"444", x"444", x"444", x"444", x"444", x"444", x"444", x"444", x"F00", x"F00"),
                                    (x"F00", x"444", x"444", x"444", x"444", x"444", x"444", x"F00", x"F00", x"F00", x"F00", x"444", x"444", x"444", x"444", x"444", x"444", x"444", x"F00", x"F00"),
                                    (x"F00", x"444", x"444", x"444", x"444", x"444", x"F00", x"F00", x"F00", x"F00", x"F00", x"F00", x"444", x"444", x"444", x"444", x"444", x"444", x"F00", x"F00"),
                                    (x"F00", x"444", x"444", x"444", x"444", x"444", x"444", x"F00", x"F00", x"F00", x"F00", x"444", x"444", x"444", x"444", x"444", x"444", x"444", x"F00", x"F00"),
                                    (x"F00", x"444", x"444", x"444", x"444", x"444", x"444", x"F00", x"F00", x"F00", x"F00", x"444", x"444", x"444", x"444", x"444", x"444", x"444", x"F00", x"F00"),
                                    (x"F00", x"444", x"444", x"444", x"444", x"444", x"444", x"F00", x"F00", x"F00", x"F00", x"444", x"444", x"444", x"444", x"444", x"444", x"444", x"F00", x"F00"),
                                    (x"F00", x"444", x"444", x"444", x"444", x"444", x"F00", x"F00", x"F00", x"F00", x"F00", x"F00", x"444", x"444", x"444", x"444", x"444", x"444", x"F00", x"F00"),
                                    (x"F00", x"444", x"444", x"444", x"444", x"444", x"444", x"F00", x"F00", x"F00", x"F00", x"444", x"444", x"444", x"444", x"444", x"444", x"444", x"F00", x"F00"),
                                    (x"F00", x"444", x"444", x"444", x"444", x"444", x"444", x"444", x"F00", x"F00", x"444", x"444", x"444", x"444", x"444", x"444", x"444", x"444", x"F00", x"F00"),
                                    (x"F00", x"444", x"444", x"444", x"444", x"444", x"444", x"444", x"F00", x"F00", x"444", x"444", x"444", x"444", x"444", x"444", x"444", x"444", x"F00", x"F00"),
                                    (x"F00", x"444", x"444", x"444", x"444", x"444", x"444", x"444", x"F00", x"F00", x"444", x"444", x"444", x"444", x"444", x"444", x"444", x"444", x"F00", x"F00"),
                                    (x"F00", x"444", x"444", x"444", x"444", x"444", x"444", x"444", x"F00", x"F00", x"444", x"444", x"444", x"444", x"444", x"444", x"444", x"444", x"F00", x"F00"),
                                    (x"F00", x"444", x"444", x"444", x"444", x"444", x"444", x"444", x"F00", x"F00", x"444", x"444", x"444", x"444", x"444", x"444", x"444", x"444", x"F00", x"F00"),
                                    (x"F00", x"444", x"444", x"444", x"444", x"444", x"444", x"F00", x"F00", x"F00", x"F00", x"444", x"444", x"444", x"444", x"444", x"444", x"444", x"F00", x"F00"),
                                    (x"F00", x"444", x"444", x"444", x"444", x"444", x"444", x"F00", x"F00", x"F00", x"F00", x"444", x"444", x"444", x"444", x"444", x"444", x"444", x"F00", x"F00"),
                                    (x"F00", x"444", x"444", x"444", x"444", x"444", x"F00", x"F00", x"F00", x"F00", x"F00", x"F00", x"444", x"444", x"444", x"444", x"444", x"444", x"F00", x"F00"),
                                    (x"F00", x"444", x"444", x"444", x"444", x"F00", x"F00", x"F00", x"F00", x"F00", x"F00", x"F00", x"F00", x"444", x"444", x"444", x"444", x"444", x"F00", x"F00"),
                                    (x"F00", x"444", x"444", x"444", x"F00", x"F00", x"F00", x"F00", x"F00", x"F00", x"F00", x"F00", x"F00", x"F00", x"444", x"444", x"444", x"444", x"F00", x"F00"),
                                    (x"F00", x"F00", x"F00", x"F00", x"F00", x"F00", x"F00", x"F00", x"F00", x"F00", x"F00", x"F00", x"F00", x"F00", x"F00", x"F00", x"F00", x"F00", x"F00", x"F00"));
    constant bishop_L : tp_cella :=((x"F00", x"F00", x"F00", x"F00", x"F00", x"F00", x"F00", x"F00", x"F00", x"F00", x"F00", x"F00", x"F00", x"F00", x"F00", x"F00", x"F00", x"F00", x"F00", x"F00"),
                                    (x"F00", x"444", x"444", x"444", x"444", x"444", x"444", x"444", x"444", x"F00", x"F00", x"444", x"444", x"444", x"444", x"444", x"444", x"444", x"F00", x"F00"),
                                    (x"F00", x"444", x"444", x"444", x"444", x"444", x"444", x"444", x"F00", x"F00", x"F00", x"F00", x"444", x"444", x"444", x"444", x"444", x"444", x"F00", x"F00"),
                                    (x"F00", x"444", x"444", x"444", x"444", x"444", x"444", x"F00", x"F00", x"F00", x"F00", x"F00", x"F00", x"444", x"444", x"444", x"444", x"444", x"F00", x"F00"),
                                    (x"F00", x"444", x"444", x"444", x"444", x"444", x"444", x"F00", x"F00", x"F00", x"F00", x"F00", x"F00", x"444", x"444", x"444", x"444", x"444", x"F00", x"F00"),
                                    (x"F00", x"444", x"444", x"444", x"444", x"444", x"444", x"F00", x"F00", x"F00", x"F00", x"F00", x"F00", x"444", x"444", x"444", x"444", x"444", x"F00", x"F00"),
                                    (x"F00", x"444", x"444", x"444", x"444", x"444", x"444", x"444", x"F00", x"F00", x"F00", x"F00", x"444", x"444", x"444", x"444", x"444", x"444", x"F00", x"F00"),
                                    (x"F00", x"444", x"444", x"444", x"444", x"444", x"444", x"444", x"444", x"F00", x"F00", x"444", x"444", x"444", x"444", x"444", x"444", x"444", x"F00", x"F00"),
                                    (x"F00", x"444", x"444", x"444", x"444", x"444", x"444", x"444", x"444", x"F00", x"F00", x"444", x"444", x"444", x"444", x"444", x"444", x"444", x"F00", x"F00"),
                                    (x"F00", x"444", x"444", x"444", x"444", x"444", x"444", x"444", x"444", x"F00", x"F00", x"444", x"444", x"444", x"444", x"444", x"444", x"444", x"F00", x"F00"),
                                    (x"F00", x"444", x"444", x"444", x"444", x"444", x"444", x"444", x"444", x"F00", x"F00", x"444", x"444", x"444", x"444", x"444", x"444", x"444", x"F00", x"F00"),
                                    (x"F00", x"444", x"444", x"444", x"444", x"444", x"444", x"444", x"444", x"F00", x"F00", x"444", x"444", x"444", x"444", x"444", x"444", x"444", x"F00", x"F00"),
                                    (x"F00", x"444", x"444", x"444", x"444", x"444", x"444", x"444", x"444", x"F00", x"F00", x"444", x"444", x"444", x"444", x"444", x"444", x"444", x"F00", x"F00"),
                                    (x"F00", x"444", x"444", x"444", x"444", x"444", x"444", x"444", x"444", x"F00", x"F00", x"444", x"444", x"444", x"444", x"444", x"444", x"444", x"F00", x"F00"),
                                    (x"F00", x"444", x"444", x"444", x"444", x"444", x"444", x"444", x"F00", x"F00", x"F00", x"F00", x"444", x"444", x"444", x"444", x"444", x"444", x"F00", x"F00"),
                                    (x"F00", x"444", x"444", x"444", x"444", x"444", x"444", x"F00", x"F00", x"F00", x"F00", x"F00", x"F00", x"444", x"444", x"444", x"444", x"444", x"F00", x"F00"),
                                    (x"F00", x"444", x"444", x"444", x"444", x"444", x"F00", x"F00", x"F00", x"F00", x"F00", x"F00", x"F00", x"F00", x"444", x"444", x"444", x"444", x"F00", x"F00"),
                                    (x"F00", x"444", x"444", x"444", x"444", x"F00", x"F00", x"F00", x"F00", x"F00", x"F00", x"F00", x"F00", x"F00", x"F00", x"444", x"444", x"444", x"F00", x"F00"),
                                    (x"F00", x"444", x"444", x"444", x"F00", x"F00", x"F00", x"F00", x"F00", x"F00", x"F00", x"F00", x"F00", x"F00", x"F00", x"F00", x"444", x"444", x"F00", x"F00"),
                                    (x"F00", x"F00", x"F00", x"F00", x"F00", x"F00", x"F00", x"F00", x"F00", x"F00", x"F00", x"F00", x"F00", x"F00", x"F00", x"F00", x"F00", x"F00", x"F00", x"F00"));
    constant tower_L : tp_cella := ((x"F00", x"F00", x"F00", x"F00", x"F00", x"F00", x"F00", x"F00", x"F00", x"F00", x"F00", x"F00", x"F00", x"F00", x"F00", x"F00", x"F00", x"F00", x"F00", x"F00"),
                                    (x"F00", x"F00", x"F00", x"F00", x"F00", x"444", x"444", x"444", x"F00", x"F00", x"F00", x"F00", x"444", x"444", x"444", x"F00", x"F00", x"F00", x"F00", x"F00"),
                                    (x"F00", x"F00", x"F00", x"F00", x"F00", x"444", x"444", x"444", x"F00", x"F00", x"F00", x"F00", x"444", x"444", x"444", x"F00", x"F00", x"F00", x"F00", x"F00"),
                                    (x"F00", x"F00", x"F00", x"F00", x"F00", x"444", x"444", x"444", x"F00", x"F00", x"F00", x"F00", x"444", x"444", x"444", x"F00", x"F00", x"F00", x"F00", x"F00"),
                                    (x"F00", x"F00", x"F00", x"F00", x"F00", x"F00", x"F00", x"F00", x"F00", x"F00", x"F00", x"F00", x"F00", x"F00", x"F00", x"F00", x"F00", x"F00", x"F00", x"F00"),
                                    (x"F00", x"F00", x"F00", x"F00", x"F00", x"F00", x"F00", x"F00", x"F00", x"F00", x"F00", x"F00", x"F00", x"F00", x"F00", x"F00", x"F00", x"F00", x"F00", x"F00"),
                                    (x"F00", x"F00", x"F00", x"F00", x"F00", x"F00", x"F00", x"F00", x"F00", x"F00", x"F00", x"F00", x"F00", x"F00", x"F00", x"F00", x"F00", x"F00", x"F00", x"F00"),
                                    (x"F00", x"F00", x"F00", x"F00", x"F00", x"F00", x"F00", x"F00", x"F00", x"F00", x"F00", x"F00", x"F00", x"F00", x"F00", x"F00", x"F00", x"F00", x"F00", x"F00"),
                                    (x"F00", x"444", x"444", x"444", x"F00", x"F00", x"F00", x"F00", x"F00", x"F00", x"F00", x"F00", x"F00", x"F00", x"F00", x"F00", x"444", x"444", x"F00", x"F00"),
                                    (x"F00", x"444", x"444", x"444", x"F00", x"F00", x"F00", x"F00", x"F00", x"F00", x"F00", x"F00", x"F00", x"F00", x"F00", x"F00", x"444", x"444", x"F00", x"F00"),
                                    (x"F00", x"444", x"444", x"444", x"F00", x"F00", x"F00", x"F00", x"F00", x"F00", x"F00", x"F00", x"F00", x"F00", x"F00", x"F00", x"444", x"444", x"F00", x"F00"),
                                    (x"F00", x"444", x"444", x"444", x"F00", x"F00", x"F00", x"F00", x"F00", x"F00", x"F00", x"F00", x"F00", x"F00", x"F00", x"F00", x"444", x"444", x"F00", x"F00"),
                                    (x"F00", x"444", x"444", x"444", x"F00", x"F00", x"F00", x"F00", x"F00", x"F00", x"F00", x"F00", x"F00", x"F00", x"F00", x"F00", x"444", x"444", x"F00", x"F00"),
                                    (x"F00", x"444", x"444", x"444", x"F00", x"F00", x"F00", x"F00", x"F00", x"F00", x"F00", x"F00", x"F00", x"F00", x"F00", x"F00", x"444", x"444", x"F00", x"F00"),
                                    (x"F00", x"444", x"444", x"444", x"F00", x"F00", x"F00", x"F00", x"F00", x"F00", x"F00", x"F00", x"F00", x"F00", x"F00", x"F00", x"444", x"444", x"F00", x"F00"),
                                    (x"F00", x"444", x"444", x"444", x"F00", x"F00", x"F00", x"F00", x"F00", x"F00", x"F00", x"F00", x"F00", x"F00", x"F00", x"F00", x"444", x"444", x"F00", x"F00"),
                                    (x"F00", x"F00", x"F00", x"F00", x"F00", x"F00", x"F00", x"F00", x"F00", x"F00", x"F00", x"F00", x"F00", x"F00", x"F00", x"F00", x"F00", x"F00", x"F00", x"F00"),
                                    (x"F00", x"F00", x"F00", x"F00", x"F00", x"F00", x"F00", x"F00", x"F00", x"F00", x"F00", x"F00", x"F00", x"F00", x"F00", x"F00", x"F00", x"F00", x"F00", x"F00"),
                                    (x"F00", x"F00", x"F00", x"F00", x"F00", x"F00", x"F00", x"F00", x"F00", x"F00", x"F00", x"F00", x"F00", x"F00", x"F00", x"F00", x"F00", x"F00", x"F00", x"F00"),
                                    (x"F00", x"F00", x"F00", x"F00", x"F00", x"F00", x"F00", x"F00", x"F00", x"F00", x"F00", x"F00", x"F00", x"F00", x"F00", x"F00", x"F00", x"F00", x"F00", x"F00"));
    constant horse_L : tp_cella := ((x"F00", x"F00", x"F00", x"F00", x"F00", x"F00", x"F00", x"F00", x"F00", x"F00", x"F00", x"F00", x"F00", x"F00", x"F00", x"F00", x"F00", x"F00", x"F00", x"F00"),
                                    (x"F00", x"444", x"444", x"444", x"444", x"444", x"444", x"444", x"F00", x"444", x"444", x"444", x"444", x"444", x"444", x"444", x"444", x"444", x"F00", x"F00"),
                                    (x"F00", x"444", x"444", x"444", x"444", x"444", x"444", x"F00", x"F00", x"F00", x"F00", x"F00", x"444", x"444", x"444", x"444", x"444", x"444", x"F00", x"F00"),
                                    (x"F00", x"444", x"444", x"444", x"444", x"444", x"F00", x"F00", x"F00", x"F00", x"F00", x"F00", x"F00", x"F00", x"F00", x"444", x"444", x"444", x"F00", x"F00"),
                                    (x"F00", x"444", x"444", x"444", x"444", x"F00", x"F00", x"F00", x"F00", x"F00", x"F00", x"F00", x"F00", x"F00", x"F00", x"444", x"444", x"444", x"F00", x"F00"),
                                    (x"F00", x"444", x"444", x"444", x"444", x"F00", x"F00", x"F00", x"F00", x"F00", x"F00", x"F00", x"F00", x"F00", x"F00", x"444", x"444", x"444", x"F00", x"F00"),
                                    (x"F00", x"444", x"444", x"444", x"444", x"F00", x"F00", x"F00", x"F00", x"F00", x"F00", x"F00", x"F00", x"F00", x"F00", x"444", x"444", x"444", x"F00", x"F00"),
                                    (x"F00", x"444", x"444", x"444", x"444", x"F00", x"F00", x"F00", x"F00", x"F00", x"F00", x"F00", x"444", x"444", x"444", x"444", x"444", x"444", x"F00", x"F00"),
                                    (x"F00", x"444", x"444", x"444", x"444", x"F00", x"F00", x"F00", x"F00", x"F00", x"F00", x"F00", x"F00", x"444", x"444", x"444", x"444", x"444", x"F00", x"F00"),
                                    (x"F00", x"444", x"444", x"444", x"444", x"F00", x"F00", x"F00", x"F00", x"F00", x"F00", x"F00", x"F00", x"F00", x"444", x"444", x"444", x"444", x"F00", x"F00"),
                                    (x"F00", x"444", x"444", x"444", x"444", x"F00", x"F00", x"F00", x"F00", x"F00", x"F00", x"F00", x"F00", x"F00", x"444", x"444", x"444", x"444", x"F00", x"F00"),
                                    (x"F00", x"444", x"444", x"444", x"444", x"F00", x"F00", x"F00", x"F00", x"F00", x"F00", x"F00", x"F00", x"F00", x"444", x"444", x"444", x"444", x"F00", x"F00"),
                                    (x"F00", x"444", x"444", x"444", x"444", x"F00", x"F00", x"F00", x"F00", x"F00", x"F00", x"F00", x"F00", x"F00", x"444", x"444", x"444", x"444", x"F00", x"F00"),
                                    (x"F00", x"444", x"444", x"444", x"444", x"F00", x"F00", x"F00", x"F00", x"F00", x"F00", x"F00", x"F00", x"444", x"444", x"444", x"444", x"444", x"F00", x"F00"),
                                    (x"F00", x"444", x"444", x"444", x"444", x"444", x"F00", x"F00", x"F00", x"F00", x"F00", x"F00", x"444", x"444", x"444", x"444", x"444", x"444", x"F00", x"F00"),
                                    (x"F00", x"444", x"444", x"444", x"444", x"444", x"444", x"F00", x"F00", x"F00", x"F00", x"444", x"444", x"444", x"444", x"444", x"444", x"444", x"F00", x"F00"),
                                    (x"F00", x"444", x"444", x"444", x"444", x"444", x"F00", x"F00", x"F00", x"F00", x"F00", x"F00", x"444", x"444", x"444", x"444", x"444", x"444", x"F00", x"F00"),
                                    (x"F00", x"444", x"444", x"444", x"444", x"F00", x"F00", x"F00", x"F00", x"F00", x"F00", x"F00", x"F00", x"444", x"444", x"444", x"444", x"444", x"F00", x"F00"),
                                    (x"F00", x"444", x"444", x"444", x"F00", x"F00", x"F00", x"F00", x"F00", x"F00", x"F00", x"F00", x"F00", x"F00", x"444", x"444", x"444", x"444", x"F00", x"F00"),
                                    (x"F00", x"F00", x"F00", x"F00", x"F00", x"F00", x"F00", x"F00", x"F00", x"F00", x"F00", x"F00", x"F00", x"F00", x"F00", x"F00", x"F00", x"F00", x"F00", x"F00"));
    -- Nero
    constant empty_D : tp_cella := ((x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000"),
                                    (x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000"),
                                    (x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000"),
                                    (x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000"),
                                    (x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000"),
                                    (x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000"),
                                    (x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000"),
                                    (x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000"),
                                    (x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000"),
                                    (x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000"),
                                    (x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000"),
                                    (x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000"),
                                    (x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000"),
                                    (x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000"),
                                    (x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000"),
                                    (x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000"),
                                    (x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000"),
                                    (x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000"),
                                    (x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000"),
                                    (x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000", x"000"));
    constant pawn_D : tp_cella :=  ((x"00F", x"00F", x"00F", x"00F", x"00F", x"00F", x"00F", x"00F", x"00F", x"00F", x"00F", x"00F", x"00F", x"00F", x"00F", x"00F", x"00F", x"00F", x"00F", x"00F"),
                                    (x"00F", x"444", x"444", x"444", x"444", x"444", x"444", x"444", x"00F", x"00F", x"00F", x"444", x"444", x"444", x"444", x"444", x"444", x"444", x"00F", x"00F"),
                                    (x"00F", x"444", x"444", x"444", x"444", x"444", x"444", x"444", x"00F", x"00F", x"00F", x"444", x"444", x"444", x"444", x"444", x"444", x"444", x"00F", x"00F"),
                                    (x"00F", x"444", x"444", x"444", x"444", x"444", x"444", x"444", x"00F", x"00F", x"00F", x"444", x"444", x"444", x"444", x"444", x"444", x"444", x"00F", x"00F"),
                                    (x"00F", x"444", x"444", x"444", x"444", x"444", x"444", x"444", x"00F", x"00F", x"00F", x"444", x"444", x"444", x"444", x"444", x"444", x"444", x"00F", x"00F"),
                                    (x"00F", x"444", x"444", x"444", x"444", x"444", x"444", x"444", x"00F", x"00F", x"00F", x"444", x"444", x"444", x"444", x"444", x"444", x"444", x"00F", x"00F"),
                                    (x"00F", x"444", x"444", x"444", x"444", x"444", x"444", x"444", x"00F", x"00F", x"00F", x"444", x"444", x"444", x"444", x"444", x"444", x"444", x"00F", x"00F"),
                                    (x"00F", x"444", x"444", x"444", x"444", x"444", x"444", x"444", x"00F", x"00F", x"00F", x"444", x"444", x"444", x"444", x"444", x"444", x"444", x"00F", x"00F"),
                                    (x"00F", x"444", x"444", x"444", x"444", x"444", x"444", x"444", x"00F", x"00F", x"00F", x"444", x"444", x"444", x"444", x"444", x"444", x"444", x"00F", x"00F"),
                                    (x"00F", x"444", x"444", x"444", x"444", x"444", x"444", x"444", x"00F", x"00F", x"00F", x"444", x"444", x"444", x"444", x"444", x"444", x"444", x"00F", x"00F"),
                                    (x"00F", x"444", x"444", x"444", x"444", x"444", x"444", x"444", x"00F", x"00F", x"00F", x"444", x"444", x"444", x"444", x"444", x"444", x"444", x"00F", x"00F"),
                                    (x"00F", x"444", x"444", x"444", x"444", x"444", x"444", x"444", x"00F", x"00F", x"00F", x"444", x"444", x"444", x"444", x"444", x"444", x"444", x"00F", x"00F"),
                                    (x"00F", x"444", x"444", x"444", x"444", x"444", x"444", x"444", x"00F", x"00F", x"00F", x"444", x"444", x"444", x"444", x"444", x"444", x"444", x"00F", x"00F"),
                                    (x"00F", x"444", x"444", x"444", x"444", x"444", x"444", x"444", x"00F", x"00F", x"00F", x"444", x"444", x"444", x"444", x"444", x"444", x"444", x"00F", x"00F"),
                                    (x"00F", x"444", x"444", x"444", x"444", x"444", x"444", x"00F", x"00F", x"00F", x"00F", x"00F", x"444", x"444", x"444", x"444", x"444", x"444", x"00F", x"00F"),
                                    (x"00F", x"444", x"444", x"444", x"444", x"444", x"444", x"00F", x"00F", x"00F", x"00F", x"00F", x"444", x"444", x"444", x"444", x"444", x"444", x"00F", x"00F"),
                                    (x"00F", x"444", x"444", x"444", x"444", x"00F", x"00F", x"00F", x"00F", x"00F", x"00F", x"00F", x"00F", x"00F", x"444", x"444", x"444", x"444", x"00F", x"00F"),
                                    (x"00F", x"444", x"444", x"444", x"00F", x"00F", x"00F", x"00F", x"00F", x"00F", x"00F", x"00F", x"00F", x"00F", x"00F", x"444", x"444", x"444", x"00F", x"00F"),
                                    (x"00F", x"444", x"444", x"00F", x"00F", x"00F", x"00F", x"00F", x"00F", x"00F", x"00F", x"00F", x"00F", x"00F", x"00F", x"00F", x"444", x"444", x"00F", x"00F"),
                                    (x"00F", x"00F", x"00F", x"00F", x"00F", x"00F", x"00F", x"00F", x"00F", x"00F", x"00F", x"00F", x"00F", x"00F", x"00F", x"00F", x"00F", x"00F", x"00F", x"00F"));
    constant king_D : tp_cella :=  ((x"00F", x"00F", x"00F", x"00F", x"00F", x"00F", x"00F", x"00F", x"00F", x"00F", x"00F", x"00F", x"00F", x"00F", x"00F", x"00F", x"00F", x"00F", x"00F", x"00F"),
                                    (x"00F", x"444", x"444", x"444", x"444", x"444", x"444", x"444", x"00F", x"00F", x"444", x"444", x"444", x"444", x"444", x"444", x"444", x"444", x"00F", x"00F"),
                                    (x"00F", x"444", x"444", x"444", x"444", x"444", x"00F", x"00F", x"00F", x"00F", x"00F", x"00F", x"444", x"444", x"444", x"444", x"444", x"444", x"00F", x"00F"),
                                    (x"00F", x"444", x"444", x"444", x"444", x"444", x"00F", x"00F", x"00F", x"00F", x"00F", x"00F", x"444", x"444", x"444", x"444", x"444", x"444", x"00F", x"00F"),
                                    (x"00F", x"444", x"444", x"444", x"444", x"444", x"444", x"444", x"00F", x"00F", x"444", x"444", x"444", x"444", x"444", x"444", x"444", x"444", x"00F", x"00F"),
                                    (x"00F", x"444", x"444", x"444", x"444", x"444", x"444", x"444", x"00F", x"00F", x"444", x"444", x"444", x"444", x"444", x"444", x"444", x"444", x"00F", x"00F"),
                                    (x"00F", x"444", x"444", x"444", x"444", x"444", x"444", x"00F", x"00F", x"00F", x"00F", x"444", x"444", x"444", x"444", x"444", x"444", x"444", x"00F", x"00F"),
                                    (x"00F", x"444", x"444", x"444", x"444", x"444", x"00F", x"00F", x"00F", x"00F", x"00F", x"00F", x"444", x"444", x"444", x"444", x"444", x"444", x"00F", x"00F"),
                                    (x"00F", x"444", x"444", x"444", x"444", x"444", x"00F", x"00F", x"00F", x"00F", x"00F", x"00F", x"444", x"444", x"444", x"444", x"444", x"444", x"00F", x"00F"),
                                    (x"00F", x"444", x"444", x"444", x"444", x"444", x"00F", x"00F", x"00F", x"00F", x"00F", x"00F", x"444", x"444", x"444", x"444", x"444", x"444", x"00F", x"00F"),
                                    (x"00F", x"444", x"444", x"444", x"444", x"00F", x"00F", x"00F", x"00F", x"00F", x"00F", x"00F", x"00F", x"444", x"444", x"444", x"444", x"444", x"00F", x"00F"),
                                    (x"00F", x"444", x"444", x"444", x"444", x"444", x"00F", x"00F", x"00F", x"00F", x"00F", x"00F", x"444", x"444", x"444", x"444", x"444", x"444", x"00F", x"00F"),
                                    (x"00F", x"444", x"444", x"444", x"444", x"444", x"444", x"00F", x"00F", x"00F", x"00F", x"444", x"444", x"444", x"444", x"444", x"444", x"444", x"00F", x"00F"),
                                    (x"00F", x"444", x"444", x"444", x"444", x"444", x"444", x"00F", x"00F", x"00F", x"00F", x"444", x"444", x"444", x"444", x"444", x"444", x"444", x"00F", x"00F"),
                                    (x"00F", x"444", x"444", x"444", x"444", x"444", x"444", x"00F", x"00F", x"00F", x"00F", x"444", x"444", x"444", x"444", x"444", x"444", x"444", x"00F", x"00F"),
                                    (x"00F", x"444", x"444", x"444", x"444", x"444", x"444", x"00F", x"00F", x"00F", x"00F", x"444", x"444", x"444", x"444", x"444", x"444", x"444", x"00F", x"00F"),
                                    (x"00F", x"444", x"444", x"444", x"444", x"444", x"00F", x"00F", x"00F", x"00F", x"00F", x"00F", x"444", x"444", x"444", x"444", x"444", x"444", x"00F", x"00F"),
                                    (x"00F", x"444", x"444", x"444", x"444", x"00F", x"00F", x"00F", x"00F", x"00F", x"00F", x"00F", x"00F", x"444", x"444", x"444", x"444", x"444", x"00F", x"00F"),
                                    (x"00F", x"444", x"444", x"444", x"00F", x"00F", x"00F", x"00F", x"00F", x"00F", x"00F", x"00F", x"00F", x"00F", x"444", x"444", x"444", x"444", x"00F", x"00F"),
                                    (x"00F", x"00F", x"00F", x"00F", x"00F", x"00F", x"00F", x"00F", x"00F", x"00F", x"00F", x"00F", x"00F", x"00F", x"00F", x"00F", x"00F", x"00F", x"00F", x"00F"));
    constant queen_D : tp_cella := ((x"00F", x"00F", x"00F", x"00F", x"00F", x"00F", x"00F", x"00F", x"00F", x"00F", x"00F", x"00F", x"00F", x"00F", x"00F", x"00F", x"00F", x"00F", x"00F", x"00F"),
                                    (x"00F", x"444", x"444", x"444", x"444", x"444", x"444", x"444", x"00F", x"00F", x"444", x"444", x"444", x"444", x"444", x"444", x"444", x"444", x"00F", x"00F"),
                                    (x"00F", x"444", x"444", x"444", x"444", x"444", x"444", x"00F", x"00F", x"00F", x"00F", x"444", x"444", x"444", x"444", x"444", x"444", x"444", x"00F", x"00F"),
                                    (x"00F", x"444", x"444", x"444", x"444", x"444", x"00F", x"00F", x"00F", x"00F", x"00F", x"00F", x"444", x"444", x"444", x"444", x"444", x"444", x"00F", x"00F"),
                                    (x"00F", x"444", x"444", x"444", x"444", x"444", x"444", x"00F", x"00F", x"00F", x"00F", x"444", x"444", x"444", x"444", x"444", x"444", x"444", x"00F", x"00F"),
                                    (x"00F", x"444", x"444", x"444", x"444", x"444", x"444", x"00F", x"00F", x"00F", x"00F", x"444", x"444", x"444", x"444", x"444", x"444", x"444", x"00F", x"00F"),
                                    (x"00F", x"444", x"444", x"444", x"444", x"444", x"444", x"00F", x"00F", x"00F", x"00F", x"444", x"444", x"444", x"444", x"444", x"444", x"444", x"00F", x"00F"),
                                    (x"00F", x"444", x"444", x"444", x"444", x"444", x"00F", x"00F", x"00F", x"00F", x"00F", x"00F", x"444", x"444", x"444", x"444", x"444", x"444", x"00F", x"00F"),
                                    (x"00F", x"444", x"444", x"444", x"444", x"444", x"444", x"00F", x"00F", x"00F", x"00F", x"444", x"444", x"444", x"444", x"444", x"444", x"444", x"00F", x"00F"),
                                    (x"00F", x"444", x"444", x"444", x"444", x"444", x"444", x"444", x"00F", x"00F", x"444", x"444", x"444", x"444", x"444", x"444", x"444", x"444", x"00F", x"00F"),
                                    (x"00F", x"444", x"444", x"444", x"444", x"444", x"444", x"444", x"00F", x"00F", x"444", x"444", x"444", x"444", x"444", x"444", x"444", x"444", x"00F", x"00F"),
                                    (x"00F", x"444", x"444", x"444", x"444", x"444", x"444", x"444", x"00F", x"00F", x"444", x"444", x"444", x"444", x"444", x"444", x"444", x"444", x"00F", x"00F"),
                                    (x"00F", x"444", x"444", x"444", x"444", x"444", x"444", x"444", x"00F", x"00F", x"444", x"444", x"444", x"444", x"444", x"444", x"444", x"444", x"00F", x"00F"),
                                    (x"00F", x"444", x"444", x"444", x"444", x"444", x"444", x"444", x"00F", x"00F", x"444", x"444", x"444", x"444", x"444", x"444", x"444", x"444", x"00F", x"00F"),
                                    (x"00F", x"444", x"444", x"444", x"444", x"444", x"444", x"00F", x"00F", x"00F", x"00F", x"444", x"444", x"444", x"444", x"444", x"444", x"444", x"00F", x"00F"),
                                    (x"00F", x"444", x"444", x"444", x"444", x"444", x"444", x"00F", x"00F", x"00F", x"00F", x"444", x"444", x"444", x"444", x"444", x"444", x"444", x"00F", x"00F"),
                                    (x"00F", x"444", x"444", x"444", x"444", x"444", x"00F", x"00F", x"00F", x"00F", x"00F", x"00F", x"444", x"444", x"444", x"444", x"444", x"444", x"00F", x"00F"),
                                    (x"00F", x"444", x"444", x"444", x"444", x"00F", x"00F", x"00F", x"00F", x"00F", x"00F", x"00F", x"00F", x"444", x"444", x"444", x"444", x"444", x"00F", x"00F"),
                                    (x"00F", x"444", x"444", x"444", x"00F", x"00F", x"00F", x"00F", x"00F", x"00F", x"00F", x"00F", x"00F", x"00F", x"444", x"444", x"444", x"444", x"00F", x"00F"),
                                    (x"00F", x"00F", x"00F", x"00F", x"00F", x"00F", x"00F", x"00F", x"00F", x"00F", x"00F", x"00F", x"00F", x"00F", x"00F", x"00F", x"00F", x"00F", x"00F", x"00F"));
    constant bishop_D : tp_cella :=((x"00F", x"00F", x"00F", x"00F", x"00F", x"00F", x"00F", x"00F", x"00F", x"00F", x"00F", x"00F", x"00F", x"00F", x"00F", x"00F", x"00F", x"00F", x"00F", x"00F"),
                                    (x"00F", x"444", x"444", x"444", x"444", x"444", x"444", x"444", x"444", x"00F", x"00F", x"444", x"444", x"444", x"444", x"444", x"444", x"444", x"00F", x"00F"),
                                    (x"00F", x"444", x"444", x"444", x"444", x"444", x"444", x"444", x"00F", x"00F", x"00F", x"00F", x"444", x"444", x"444", x"444", x"444", x"444", x"00F", x"00F"),
                                    (x"00F", x"444", x"444", x"444", x"444", x"444", x"444", x"00F", x"00F", x"00F", x"00F", x"00F", x"00F", x"444", x"444", x"444", x"444", x"444", x"00F", x"00F"),
                                    (x"00F", x"444", x"444", x"444", x"444", x"444", x"444", x"00F", x"00F", x"00F", x"00F", x"00F", x"00F", x"444", x"444", x"444", x"444", x"444", x"00F", x"00F"),
                                    (x"00F", x"444", x"444", x"444", x"444", x"444", x"444", x"00F", x"00F", x"00F", x"00F", x"00F", x"00F", x"444", x"444", x"444", x"444", x"444", x"00F", x"00F"),
                                    (x"00F", x"444", x"444", x"444", x"444", x"444", x"444", x"444", x"00F", x"00F", x"00F", x"00F", x"444", x"444", x"444", x"444", x"444", x"444", x"00F", x"00F"),
                                    (x"00F", x"444", x"444", x"444", x"444", x"444", x"444", x"444", x"444", x"00F", x"00F", x"444", x"444", x"444", x"444", x"444", x"444", x"444", x"00F", x"00F"),
                                    (x"00F", x"444", x"444", x"444", x"444", x"444", x"444", x"444", x"444", x"00F", x"00F", x"444", x"444", x"444", x"444", x"444", x"444", x"444", x"00F", x"00F"),
                                    (x"00F", x"444", x"444", x"444", x"444", x"444", x"444", x"444", x"444", x"00F", x"00F", x"444", x"444", x"444", x"444", x"444", x"444", x"444", x"00F", x"00F"),
                                    (x"00F", x"444", x"444", x"444", x"444", x"444", x"444", x"444", x"444", x"00F", x"00F", x"444", x"444", x"444", x"444", x"444", x"444", x"444", x"00F", x"00F"),
                                    (x"00F", x"444", x"444", x"444", x"444", x"444", x"444", x"444", x"444", x"00F", x"00F", x"444", x"444", x"444", x"444", x"444", x"444", x"444", x"00F", x"00F"),
                                    (x"00F", x"444", x"444", x"444", x"444", x"444", x"444", x"444", x"444", x"00F", x"00F", x"444", x"444", x"444", x"444", x"444", x"444", x"444", x"00F", x"00F"),
                                    (x"00F", x"444", x"444", x"444", x"444", x"444", x"444", x"444", x"444", x"00F", x"00F", x"444", x"444", x"444", x"444", x"444", x"444", x"444", x"00F", x"00F"),
                                    (x"00F", x"444", x"444", x"444", x"444", x"444", x"444", x"444", x"00F", x"00F", x"00F", x"00F", x"444", x"444", x"444", x"444", x"444", x"444", x"00F", x"00F"),
                                    (x"00F", x"444", x"444", x"444", x"444", x"444", x"444", x"00F", x"00F", x"00F", x"00F", x"00F", x"00F", x"444", x"444", x"444", x"444", x"444", x"00F", x"00F"),
                                    (x"00F", x"444", x"444", x"444", x"444", x"444", x"00F", x"00F", x"00F", x"00F", x"00F", x"00F", x"00F", x"00F", x"444", x"444", x"444", x"444", x"00F", x"00F"),
                                    (x"00F", x"444", x"444", x"444", x"444", x"00F", x"00F", x"00F", x"00F", x"00F", x"00F", x"00F", x"00F", x"00F", x"00F", x"444", x"444", x"444", x"00F", x"00F"),
                                    (x"00F", x"444", x"444", x"444", x"00F", x"00F", x"00F", x"00F", x"00F", x"00F", x"00F", x"00F", x"00F", x"00F", x"00F", x"00F", x"444", x"444", x"00F", x"00F"),
                                    (x"00F", x"00F", x"00F", x"00F", x"00F", x"00F", x"00F", x"00F", x"00F", x"00F", x"00F", x"00F", x"00F", x"00F", x"00F", x"00F", x"00F", x"00F", x"00F", x"00F"));
    constant tower_D : tp_cella := ((x"00F", x"00F", x"00F", x"00F", x"00F", x"00F", x"00F", x"00F", x"00F", x"00F", x"00F", x"00F", x"00F", x"00F", x"00F", x"00F", x"00F", x"00F", x"00F", x"00F"),
                                    (x"00F", x"00F", x"00F", x"00F", x"00F", x"444", x"444", x"444", x"00F", x"00F", x"00F", x"00F", x"444", x"444", x"444", x"00F", x"00F", x"00F", x"00F", x"00F"),
                                    (x"00F", x"00F", x"00F", x"00F", x"00F", x"444", x"444", x"444", x"00F", x"00F", x"00F", x"00F", x"444", x"444", x"444", x"00F", x"00F", x"00F", x"00F", x"00F"),
                                    (x"00F", x"00F", x"00F", x"00F", x"00F", x"444", x"444", x"444", x"00F", x"00F", x"00F", x"00F", x"444", x"444", x"444", x"00F", x"00F", x"00F", x"00F", x"00F"),
                                    (x"00F", x"00F", x"00F", x"00F", x"00F", x"00F", x"00F", x"00F", x"00F", x"00F", x"00F", x"00F", x"00F", x"00F", x"00F", x"00F", x"00F", x"00F", x"00F", x"00F"),
                                    (x"00F", x"00F", x"00F", x"00F", x"00F", x"00F", x"00F", x"00F", x"00F", x"00F", x"00F", x"00F", x"00F", x"00F", x"00F", x"00F", x"00F", x"00F", x"00F", x"00F"),
                                    (x"00F", x"00F", x"00F", x"00F", x"00F", x"00F", x"00F", x"00F", x"00F", x"00F", x"00F", x"00F", x"00F", x"00F", x"00F", x"00F", x"00F", x"00F", x"00F", x"00F"),
                                    (x"00F", x"00F", x"00F", x"00F", x"00F", x"00F", x"00F", x"00F", x"00F", x"00F", x"00F", x"00F", x"00F", x"00F", x"00F", x"00F", x"00F", x"00F", x"00F", x"00F"),
                                    (x"00F", x"444", x"444", x"444", x"00F", x"00F", x"00F", x"00F", x"00F", x"00F", x"00F", x"00F", x"00F", x"00F", x"00F", x"00F", x"444", x"444", x"00F", x"00F"),
                                    (x"00F", x"444", x"444", x"444", x"00F", x"00F", x"00F", x"00F", x"00F", x"00F", x"00F", x"00F", x"00F", x"00F", x"00F", x"00F", x"444", x"444", x"00F", x"00F"),
                                    (x"00F", x"444", x"444", x"444", x"00F", x"00F", x"00F", x"00F", x"00F", x"00F", x"00F", x"00F", x"00F", x"00F", x"00F", x"00F", x"444", x"444", x"00F", x"00F"),
                                    (x"00F", x"444", x"444", x"444", x"00F", x"00F", x"00F", x"00F", x"00F", x"00F", x"00F", x"00F", x"00F", x"00F", x"00F", x"00F", x"444", x"444", x"00F", x"00F"),
                                    (x"00F", x"444", x"444", x"444", x"00F", x"00F", x"00F", x"00F", x"00F", x"00F", x"00F", x"00F", x"00F", x"00F", x"00F", x"00F", x"444", x"444", x"00F", x"00F"),
                                    (x"00F", x"444", x"444", x"444", x"00F", x"00F", x"00F", x"00F", x"00F", x"00F", x"00F", x"00F", x"00F", x"00F", x"00F", x"00F", x"444", x"444", x"00F", x"00F"),
                                    (x"00F", x"444", x"444", x"444", x"00F", x"00F", x"00F", x"00F", x"00F", x"00F", x"00F", x"00F", x"00F", x"00F", x"00F", x"00F", x"444", x"444", x"00F", x"00F"),
                                    (x"00F", x"444", x"444", x"444", x"00F", x"00F", x"00F", x"00F", x"00F", x"00F", x"00F", x"00F", x"00F", x"00F", x"00F", x"00F", x"444", x"444", x"00F", x"00F"),
                                    (x"00F", x"00F", x"00F", x"00F", x"00F", x"00F", x"00F", x"00F", x"00F", x"00F", x"00F", x"00F", x"00F", x"00F", x"00F", x"00F", x"00F", x"00F", x"00F", x"00F"),
                                    (x"00F", x"00F", x"00F", x"00F", x"00F", x"00F", x"00F", x"00F", x"00F", x"00F", x"00F", x"00F", x"00F", x"00F", x"00F", x"00F", x"00F", x"00F", x"00F", x"00F"),
                                    (x"00F", x"00F", x"00F", x"00F", x"00F", x"00F", x"00F", x"00F", x"00F", x"00F", x"00F", x"00F", x"00F", x"00F", x"00F", x"00F", x"00F", x"00F", x"00F", x"00F"),
                                    (x"00F", x"00F", x"00F", x"00F", x"00F", x"00F", x"00F", x"00F", x"00F", x"00F", x"00F", x"00F", x"00F", x"00F", x"00F", x"00F", x"00F", x"00F", x"00F", x"00F"));
    constant horse_D : tp_cella := ((x"00F", x"00F", x"00F", x"00F", x"00F", x"00F", x"00F", x"00F", x"00F", x"00F", x"00F", x"00F", x"00F", x"00F", x"00F", x"00F", x"00F", x"00F", x"00F", x"00F"),
                                    (x"00F", x"444", x"444", x"444", x"444", x"444", x"444", x"444", x"00F", x"444", x"444", x"444", x"444", x"444", x"444", x"444", x"444", x"444", x"00F", x"00F"),
                                    (x"00F", x"444", x"444", x"444", x"444", x"444", x"444", x"00F", x"00F", x"00F", x"00F", x"00F", x"444", x"444", x"444", x"444", x"444", x"444", x"00F", x"00F"),
                                    (x"00F", x"444", x"444", x"444", x"444", x"444", x"00F", x"00F", x"00F", x"00F", x"00F", x"00F", x"00F", x"00F", x"00F", x"444", x"444", x"444", x"00F", x"00F"),
                                    (x"00F", x"444", x"444", x"444", x"444", x"00F", x"00F", x"00F", x"00F", x"00F", x"00F", x"00F", x"00F", x"00F", x"00F", x"444", x"444", x"444", x"00F", x"00F"),
                                    (x"00F", x"444", x"444", x"444", x"444", x"00F", x"00F", x"00F", x"00F", x"00F", x"00F", x"00F", x"00F", x"00F", x"00F", x"444", x"444", x"444", x"00F", x"00F"),
                                    (x"00F", x"444", x"444", x"444", x"444", x"00F", x"00F", x"00F", x"00F", x"00F", x"00F", x"00F", x"00F", x"00F", x"00F", x"444", x"444", x"444", x"00F", x"00F"),
                                    (x"00F", x"444", x"444", x"444", x"444", x"00F", x"00F", x"00F", x"00F", x"00F", x"00F", x"00F", x"444", x"444", x"444", x"444", x"444", x"444", x"00F", x"00F"),
                                    (x"00F", x"444", x"444", x"444", x"444", x"00F", x"00F", x"00F", x"00F", x"00F", x"00F", x"00F", x"00F", x"444", x"444", x"444", x"444", x"444", x"00F", x"00F"),
                                    (x"00F", x"444", x"444", x"444", x"444", x"00F", x"00F", x"00F", x"00F", x"00F", x"00F", x"00F", x"00F", x"00F", x"444", x"444", x"444", x"444", x"00F", x"00F"),
                                    (x"00F", x"444", x"444", x"444", x"444", x"00F", x"00F", x"00F", x"00F", x"00F", x"00F", x"00F", x"00F", x"00F", x"444", x"444", x"444", x"444", x"00F", x"00F"),
                                    (x"00F", x"444", x"444", x"444", x"444", x"00F", x"00F", x"00F", x"00F", x"00F", x"00F", x"00F", x"00F", x"00F", x"444", x"444", x"444", x"444", x"00F", x"00F"),
                                    (x"00F", x"444", x"444", x"444", x"444", x"00F", x"00F", x"00F", x"00F", x"00F", x"00F", x"00F", x"00F", x"00F", x"444", x"444", x"444", x"444", x"00F", x"00F"),
                                    (x"00F", x"444", x"444", x"444", x"444", x"00F", x"00F", x"00F", x"00F", x"00F", x"00F", x"00F", x"00F", x"444", x"444", x"444", x"444", x"444", x"00F", x"00F"),
                                    (x"00F", x"444", x"444", x"444", x"444", x"444", x"00F", x"00F", x"00F", x"00F", x"00F", x"00F", x"444", x"444", x"444", x"444", x"444", x"444", x"00F", x"00F"),
                                    (x"00F", x"444", x"444", x"444", x"444", x"444", x"444", x"00F", x"00F", x"00F", x"00F", x"444", x"444", x"444", x"444", x"444", x"444", x"444", x"00F", x"00F"),
                                    (x"00F", x"444", x"444", x"444", x"444", x"444", x"00F", x"00F", x"00F", x"00F", x"00F", x"00F", x"444", x"444", x"444", x"444", x"444", x"444", x"00F", x"00F"),
                                    (x"00F", x"444", x"444", x"444", x"444", x"00F", x"00F", x"00F", x"00F", x"00F", x"00F", x"00F", x"00F", x"444", x"444", x"444", x"444", x"444", x"00F", x"00F"),
                                    (x"00F", x"444", x"444", x"444", x"00F", x"00F", x"00F", x"00F", x"00F", x"00F", x"00F", x"00F", x"00F", x"00F", x"444", x"444", x"444", x"444", x"00F", x"00F"),
                                    (x"00F", x"00F", x"00F", x"00F", x"00F", x"00F", x"00F", x"00F", x"00F", x"00F", x"00F", x"00F", x"00F", x"00F", x"00F", x"00F", x"00F", x"00F", x"00F", x"00F"));
---------------------------------------------------------------------------------------------------------------------------------
-- SIGNAL DECLARATION                                                                                                      
--------------------------------------------------------------------------------------------------------------------------------- 
    signal si_curs_x_reg0:  integer range 0 to 8        := 0                ;
    signal si_curs_y_reg0:  integer range 0 to 8        := 0                ;   
    signal si_curs_x_reg1:  integer range 0 to 8        := 0                ;
    signal si_curs_y_reg1:  integer range 0 to 8        := 0                ; 
    signal si_curs_x     :  integer range 0 to 8        := 0                ;
    signal si_curs_y     :  integer range 0 to 8        := 0                ;
    signal st_stato      :  tp_stato                    := IDLE             ;
    signal st_stato_dopo :  tp_stato                    := IDLE             ;
    signal sv_delay_ms   :  std_logic_vector(11 downto 0):= (others => '0') ;
    signal ss_delay_en   :  std_logic                   := '0'              ;
    signal ss_delay_done :  std_logic                   := '0'              ;
    signal ss_lamp_on    :  std_logic                   := '0'              ;
    signal st_cursore    :  tp_cella                    := empty_L          ;
    signal st_lamp_on    :  tp_cella                    := empty_L          ;
    signal st_lamp_off   :  tp_cella                    := empty_L          ;
    signal st_lamp_off1  :  tp_cella                    := empty_L          ;

    signal clk_div       :  unsigned(1 downto 0)        := (others => '0')  ;
    signal sv_r          :  std_logic_vector(3 downto 0):= "0111"           ;
    signal sv_b          :  std_logic_vector(3 downto 0):= "0111"           ;
    signal sv_g          :  std_logic_vector(3 downto 0):= "0111"           ;
    signal sv_v_cnt      :  unsigned(10 downto 0)       := (others => '0')  ;
    signal sv_h_cnt      :  unsigned(10 downto 0)       := (others => '0')  ;
    signal ss_ack        :  std_logic                   := '0'              ;
    signal sv_numero     :  std_logic_vector(5 downto 0):= "000000"         ;
    signal sv_tipo       :  std_logic_vector(3 downto 0):= "0000"           ;
    signal sv_x_matrix   :  unsigned(10 downto 0)       := (others => '0')  ;
    signal sv_y_matrix   :  unsigned(10 downto 0)       := (others => '0')  ;    
    --scacchiera 
    --A0 A1 A2 A3 A4 A5 A6 A7
    --B0 B1 B2 B3 B4 B5 B6 B7
    --C0 C1 C2 C3 C4 C5 C6 C7
    --D0 D1 D2 D3 D4 D5 D6 D7
    --E0 E1 E2 E3 E4 E5 E6 E7
    --F0 F1 F2 F3 F4 F5 F6 F7
    --G0 G1 G2 G3 G4 G5 G6 G7
    --H0 H1 H2 H3 H4 H5 H6 H7
    signal A0, A1, A2, A3, A4, A5, A6, A7   :   tp_cella := empty_L;
    signal B0, B1, B2, B3, B4, B5, B6, B7   :   tp_cella := empty_L;
    signal C0, C1, C2, C3, C4, C5, C6, C7   :   tp_cella := empty_L;
    signal D0, D1, D2, D3, D4, D5, D6, D7   :   tp_cella := empty_L;
    signal E0, E1, E2, E3, E4, E5, E6, E7   :   tp_cella := empty_L;
    signal F0, F1, F2, F3, F4, F5, F6, F7   :   tp_cella := empty_L;
    signal G0, G1, G2, G3, G4, G5, G6, G7   :   tp_cella := empty_L;
    signal H0, H1, H2, H3, H4, H5, H6, H7   :   tp_cella := empty_L;
    
    begin
---------------------------------------------------------------------------------------------------------------------------------
-- ASSEGNAZIONE SEGNALI IN                                                                                                            
---------------------------------------------------------------------------------------------------------------------------------    
        sv_v_cnt        <= unsigned(FRM_i_V_CNT) ;
        sv_h_cnt        <= unsigned(FRM_i_H_CNT) ;
        si_curs_x_reg0  <= to_integer(unsigned(FRM_i_CURS_X));
        si_curs_y_reg0  <= to_integer(unsigned(FRM_i_CURS_Y));
        ss_delay_done   <= FRM_i_DONE            ;
---------------------------------------------------------------------------------------------------------------------------------
-- ASSEGNAZIONE SEGNALI OUT                                                                                                            
---------------------------------------------------------------------------------------------------------------------------------
        FRM_o_ACK       <= ss_ack     ;
        FRM_o_DELAY_MS  <= sv_delay_ms;
        FRM_o_DELAY_EN  <= ss_delay_en;

        RICREAZIONE_SCACCHIERA: process (FRM_i_CLK_100M) begin
            if (rising_edge(FRM_i_CLK_100M)) then
                clk_div <= clk_div + 1;
                ss_ack <= '0';
                if(clk_div = 3) then
                    clk_div <= (others => '0');
                    ss_ack <= '1';
                if(ss_ack <= '1') then
                    -- Divido numero e tipologia di PEZZO
                    sv_numero   <=  FRM_i_PIECE(9 downto 4);
                    sv_tipo     <=  FRM_i_PIECE(3 downto 0);
                    
                    case sv_numero is 
                        when "000000" => -- A0 / casella : 0
                            case sv_tipo is
                                when "0000" => A0 <= empty_L ; -- vuoto bianco
                                when "0001" => A0 <= pawn_L  ; -- pedone bianco
                                when "0010" => A0 <= king_L  ; -- re bianco
                                when "0011" => A0 <= queen_L ; -- regina bianco
                                when "0100" => A0 <= bishop_L; -- alfiere bianco
                                when "0101" => A0 <= tower_L ; -- torre bianco
                                when "0110" => A0 <= horse_L ; -- cavallo bianco
                                when "1000" => A0 <= empty_D ; -- vuoto bianco  
                                when "1001" => A0 <= pawn_D  ; -- pedone nero 
                                when "1010" => A0 <= king_D  ; -- re nero     
                                when "1011" => A0 <= queen_D ; -- regina nero 
                                when "1100" => A0 <= bishop_D; -- alfiere nero
                                when "1101" => A0 <= tower_D ; -- torre nero  
                                when "1110" => A0 <= horse_D ; -- cavallo nero
                                when others => A0 <= empty_L ; -- vuoto bianco default
                            end case;
                        when "000001" => -- A1 / casella : 1
                            case sv_tipo is
                                when "0000" => A1 <= empty_L ; -- vuoto bianco
                                when "0001" => A1 <= pawn_L  ; -- pedone bianco
                                when "0010" => A1 <= king_L  ; -- re bianco
                                when "0011" => A1 <= queen_L ; -- regina bianco
                                when "0100" => A1 <= bishop_L; -- alfiere bianco
                                when "0101" => A1 <= tower_L ; -- torre bianco
                                when "0110" => A1 <= horse_L ; -- cavallo bianco
                                when "1000" => A1 <= empty_D ; -- vuoto bianco  
                                when "1001" => A1 <= pawn_D  ; -- pedone nero 
                                when "1010" => A1 <= king_D  ; -- re nero     
                                when "1011" => A1 <= queen_D ; -- regina nero 
                                when "1100" => A1 <= bishop_D; -- alfiere nero
                                when "1101" => A1 <= tower_D ; -- torre nero  
                                when "1110" => A1 <= horse_D ; -- cavallo nero
                                when others => A1 <= empty_L ; -- vuoto bianco default
                            end case;
                        when "000010" => -- A2 / casella : 2
                            case sv_tipo is
                                when "0000" => A2 <= empty_L ; -- vuoto bianco
                                when "0001" => A2 <= pawn_L  ; -- pedone bianco
                                when "0010" => A2 <= king_L  ; -- re bianco
                                when "0011" => A2 <= queen_L ; -- regina bianco
                                when "0100" => A2 <= bishop_L; -- alfiere bianco
                                when "0101" => A2 <= tower_L ; -- torre bianco
                                when "0110" => A2 <= horse_L ; -- cavallo bianco
                                when "1000" => A2 <= empty_D ; -- vuoto bianco  
                                when "1001" => A2 <= pawn_D  ; -- pedone nero 
                                when "1010" => A2 <= king_D  ; -- re nero     
                                when "1011" => A2 <= queen_D ; -- regina nero 
                                when "1100" => A2 <= bishop_D; -- alfiere nero
                                when "1101" => A2 <= tower_D ; -- torre nero  
                                when "1110" => A2 <= horse_D ; -- cavallo nero
                                when others => A2 <= empty_L ; -- vuoto bianco default
                            end case;
                        when "000011" => -- A3 / casella : 3
                            case sv_tipo is
                                when "0000" => A3 <= empty_L ; -- vuoto bianco
                                when "0001" => A3 <= pawn_L  ; -- pedone bianco
                                when "0010" => A3 <= king_L  ; -- re bianco
                                when "0011" => A3 <= queen_L ; -- regina bianco
                                when "0100" => A3 <= bishop_L; -- alfiere bianco
                                when "0101" => A3 <= tower_L ; -- torre bianco
                                when "0110" => A3 <= horse_L ; -- cavallo bianco
                                when "1000" => A3 <= empty_D ; -- vuoto bianco  
                                when "1001" => A3 <= pawn_D  ; -- pedone nero 
                                when "1010" => A3 <= king_D  ; -- re nero     
                                when "1011" => A3 <= queen_D ; -- regina nero 
                                when "1100" => A3 <= bishop_D; -- alfiere nero
                                when "1101" => A3 <= tower_D ; -- torre nero  
                                when "1110" => A3 <= horse_D ; -- cavallo nero
                                when others => A3 <= empty_L ; -- vuoto bianco default
                            end case;
                        when "000100" => -- A4 / casella : 4
                            case sv_tipo is
                                when "0000" => A4 <= empty_L ; -- vuoto bianco
                                when "0001" => A4 <= pawn_L  ; -- pedone bianco
                                when "0010" => A4 <= king_L  ; -- re bianco
                                when "0011" => A4 <= queen_L ; -- regina bianco
                                when "0100" => A4 <= bishop_L; -- alfiere bianco
                                when "0101" => A4 <= tower_L ; -- torre bianco
                                when "0110" => A4 <= horse_L ; -- cavallo bianco
                                when "1000" => A4 <= empty_D ; -- vuoto bianco  
                                when "1001" => A4 <= pawn_D  ; -- pedone nero 
                                when "1010" => A4 <= king_D  ; -- re nero     
                                when "1011" => A4 <= queen_D ; -- regina nero 
                                when "1100" => A4 <= bishop_D; -- alfiere nero
                                when "1101" => A4 <= tower_D ; -- torre nero  
                                when "1110" => A4 <= horse_D ; -- cavallo nero
                                when others => A4 <= empty_L ; -- vuoto bianco default
                            end case;
                        when "000101" => -- A5 / casella : 5
                            case sv_tipo is
                                when "0000" => A5 <= empty_L ; -- vuoto bianco
                                when "0001" => A5 <= pawn_L  ; -- pedone bianco
                                when "0010" => A5 <= king_L  ; -- re bianco
                                when "0011" => A5 <= queen_L ; -- regina bianco
                                when "0100" => A5 <= bishop_L; -- alfiere bianco
                                when "0101" => A5 <= tower_L ; -- torre bianco
                                when "0110" => A5 <= horse_L ; -- cavallo bianco
                                when "1000" => A5 <= empty_D ; -- vuoto bianco  
                                when "1001" => A5 <= pawn_D  ; -- pedone nero 
                                when "1010" => A5 <= king_D  ; -- re nero     
                                when "1011" => A5 <= queen_D ; -- regina nero 
                                when "1100" => A5 <= bishop_D; -- alfiere nero
                                when "1101" => A5 <= tower_D ; -- torre nero  
                                when "1110" => A5 <= horse_D ; -- cavallo nero
                                when others => A5 <= empty_L ; -- vuoto bianco default
                            end case;
                        when "000110" => -- A6 / casella : 6
                            case sv_tipo is
                                when "0000" => A6 <= empty_L ; -- vuoto bianco
                                when "0001" => A6 <= pawn_L  ; -- pedone bianco
                                when "0010" => A6 <= king_L  ; -- re bianco
                                when "0011" => A6 <= queen_L ; -- regina bianco
                                when "0100" => A6 <= bishop_L; -- alfiere bianco
                                when "0101" => A6 <= tower_L ; -- torre bianco
                                when "0110" => A6 <= horse_L ; -- cavallo bianco
                                when "1000" => A6 <= empty_D ; -- vuoto bianco  
                                when "1001" => A6 <= pawn_D  ; -- pedone nero 
                                when "1010" => A6 <= king_D  ; -- re nero     
                                when "1011" => A6 <= queen_D ; -- regina nero 
                                when "1100" => A6 <= bishop_D; -- alfiere nero
                                when "1101" => A6 <= tower_D ; -- torre nero  
                                when "1110" => A6 <= horse_D ; -- cavallo nero
                                when others => A6 <= empty_L ; -- vuoto bianco default
                            end case;
                        when "000111" => -- A7 / casella : 7
                            case sv_tipo is
                                when "0000" => A7 <= empty_L ; -- vuoto bianco
                                when "0001" => A7 <= pawn_L  ; -- pedone bianco
                                when "0010" => A7 <= king_L  ; -- re bianco
                                when "0011" => A7 <= queen_L ; -- regina bianco
                                when "0100" => A7 <= bishop_L; -- alfiere bianco
                                when "0101" => A7 <= tower_L ; -- torre bianco
                                when "0110" => A7 <= horse_L ; -- cavallo bianco
                                when "1000" => A7 <= empty_D ; -- vuoto bianco  
                                when "1001" => A7 <= pawn_D  ; -- pedone nero 
                                when "1010" => A7 <= king_D  ; -- re nero     
                                when "1011" => A7 <= queen_D ; -- regina nero 
                                when "1100" => A7 <= bishop_D; -- alfiere nero
                                when "1101" => A7 <= tower_D ; -- torre nero  
                                when "1110" => A7 <= horse_D ; -- cavallo nero
                                when others => A7 <= empty_L ; -- vuoto bianco default
                            end case;
                        when "001000" => -- B0 / casella : 8
                            case sv_tipo is
                                when "0000" => B0 <= empty_L ; -- vuoto bianco
                                when "0001" => B0 <= pawn_L  ; -- pedone bianco
                                when "0010" => B0 <= king_L  ; -- re bianco
                                when "0011" => B0 <= queen_L ; -- regina bianco
                                when "0100" => B0 <= bishop_L; -- alfiere bianco
                                when "0101" => B0 <= tower_L ; -- torre bianco
                                when "0110" => B0 <= horse_L ; -- cavallo bianco
                                when "1000" => B0 <= empty_D ; -- vuoto bianco  
                                when "1001" => B0 <= pawn_D  ; -- pedone nero 
                                when "1010" => B0 <= king_D  ; -- re nero     
                                when "1011" => B0 <= queen_D ; -- regina nero 
                                when "1100" => B0 <= bishop_D; -- alfiere nero
                                when "1101" => B0 <= tower_D ; -- torre nero  
                                when "1110" => B0 <= horse_D ; -- cavallo nero
                                when others => B0 <= empty_L ; -- vuoto bianco default
                            end case;
                        when "001001" => -- B1 / casella : 9 
                            case sv_tipo is
                                when "0000" => B1 <= empty_L ; -- vuoto bianco
                                when "0001" => B1 <= pawn_L  ; -- pedone bianco
                                when "0010" => B1 <= king_L  ; -- re bianco
                                when "0011" => B1 <= queen_L ; -- regina bianco
                                when "0100" => B1 <= bishop_L; -- alfiere bianco
                                when "0101" => B1 <= tower_L ; -- torre bianco
                                when "0110" => B1 <= horse_L ; -- cavallo bianco
                                when "1000" => B1 <= empty_D ; -- vuoto bianco  
                                when "1001" => B1 <= pawn_D  ; -- pedone nero 
                                when "1010" => B1 <= king_D  ; -- re nero     
                                when "1011" => B1 <= queen_D ; -- regina nero 
                                when "1100" => B1 <= bishop_D; -- alfiere nero
                                when "1101" => B1 <= tower_D ; -- torre nero  
                                when "1110" => B1 <= horse_D ; -- cavallo nero
                                when others => B1 <= empty_L ; -- vuoto bianco default
                            end case;
                        when "001010" => -- B2 / casella : 10
                            case sv_tipo is
                                when "0000" => B2 <= empty_L ; -- vuoto bianco
                                when "0001" => B2 <= pawn_L  ; -- pedone bianco
                                when "0010" => B2 <= king_L  ; -- re bianco
                                when "0011" => B2 <= queen_L ; -- regina bianco
                                when "0100" => B2 <= bishop_L; -- alfiere bianco
                                when "0101" => B2 <= tower_L ; -- torre bianco
                                when "0110" => B2 <= horse_L ; -- cavallo bianco
                                when "1000" => B2 <= empty_D ; -- vuoto bianco  
                                when "1001" => B2 <= pawn_D  ; -- pedone nero 
                                when "1010" => B2 <= king_D  ; -- re nero     
                                when "1011" => B2 <= queen_D ; -- regina nero 
                                when "1100" => B2 <= bishop_D; -- alfiere nero
                                when "1101" => B2 <= tower_D ; -- torre nero  
                                when "1110" => B2 <= horse_D ; -- cavallo nero
                                when others => B2 <= empty_L ; -- vuoto bianco default
                            end case;
                        when "001011" => -- B3 / casella : 11
                            case sv_tipo is
                                when "0000" => B3 <= empty_L ; -- vuoto bianco
                                when "0001" => B3 <= pawn_L  ; -- pedone bianco
                                when "0010" => B3 <= king_L  ; -- re bianco
                                when "0011" => B3 <= queen_L ; -- regina bianco
                                when "0100" => B3 <= bishop_L; -- alfiere bianco
                                when "0101" => B3 <= tower_L ; -- torre bianco
                                when "0110" => B3 <= horse_L ; -- cavallo bianco
                                when "1000" => B3 <= empty_D ; -- vuoto bianco  
                                when "1001" => B3 <= pawn_D  ; -- pedone nero 
                                when "1010" => B3 <= king_D  ; -- re nero     
                                when "1011" => B3 <= queen_D ; -- regina nero 
                                when "1100" => B3 <= bishop_D; -- alfiere nero
                                when "1101" => B3 <= tower_D ; -- torre nero  
                                when "1110" => B3 <= horse_D ; -- cavallo nero
                                when others => B3 <= empty_L ; -- vuoto bianco default
                            end case;
                        when "001100" => -- B4 / casella : 12
                            case sv_tipo is
                                when "0000" => B4 <= empty_L ; -- vuoto bianco
                                when "0001" => B4 <= pawn_L  ; -- pedone bianco
                                when "0010" => B4 <= king_L  ; -- re bianco
                                when "0011" => B4 <= queen_L ; -- regina bianco
                                when "0100" => B4 <= bishop_L; -- alfiere bianco
                                when "0101" => B4 <= tower_L ; -- torre bianco
                                when "0110" => B4 <= horse_L ; -- cavallo bianco
                                when "1000" => B4 <= empty_D ; -- vuoto bianco  
                                when "1001" => B4 <= pawn_D  ; -- pedone nero 
                                when "1010" => B4 <= king_D  ; -- re nero     
                                when "1011" => B4 <= queen_D ; -- regina nero 
                                when "1100" => B4 <= bishop_D; -- alfiere nero
                                when "1101" => B4 <= tower_D ; -- torre nero  
                                when "1110" => B4 <= horse_D ; -- cavallo nero
                                when others => B4 <= empty_L ; -- vuoto bianco default
                            end case;
                        when "001101" => -- B5 / casella : 13
                            case sv_tipo is
                                when "0000" => B5 <= empty_L ; -- vuoto bianco
                                when "0001" => B5 <= pawn_L  ; -- pedone bianco
                                when "0010" => B5 <= king_L  ; -- re bianco
                                when "0011" => B5 <= queen_L ; -- regina bianco
                                when "0100" => B5 <= bishop_L; -- alfiere bianco
                                when "0101" => B5 <= tower_L ; -- torre bianco
                                when "0110" => B5 <= horse_L ; -- cavallo bianco
                                when "1000" => B5 <= empty_D ; -- vuoto bianco  
                                when "1001" => B5 <= pawn_D  ; -- pedone nero 
                                when "1010" => B5 <= king_D  ; -- re nero     
                                when "1011" => B5 <= queen_D ; -- regina nero 
                                when "1100" => B5 <= bishop_D; -- alfiere nero
                                when "1101" => B5 <= tower_D ; -- torre nero  
                                when "1110" => B5 <= horse_D ; -- cavallo nero
                                when others => B5 <= empty_L ; -- vuoto bianco default
                            end case;
                        when "001110" => -- B6 / casella : 14
                            case sv_tipo is
                                when "0000" => B6 <= empty_L ; -- vuoto bianco
                                when "0001" => B6 <= pawn_L  ; -- pedone bianco
                                when "0010" => B6 <= king_L  ; -- re bianco
                                when "0011" => B6 <= queen_L ; -- regina bianco
                                when "0100" => B6 <= bishop_L; -- alfiere bianco
                                when "0101" => B6 <= tower_L ; -- torre bianco
                                when "0110" => B6 <= horse_L ; -- cavallo bianco
                                when "1000" => B6 <= empty_D ; -- vuoto bianco  
                                when "1001" => B6 <= pawn_D  ; -- pedone nero 
                                when "1010" => B6 <= king_D  ; -- re nero     
                                when "1011" => B6 <= queen_D ; -- regina nero 
                                when "1100" => B6 <= bishop_D; -- alfiere nero
                                when "1101" => B6 <= tower_D ; -- torre nero  
                                when "1110" => B6 <= horse_D ; -- cavallo nero
                                when others => B6 <= empty_L ; -- vuoto bianco default
                            end case;
                        when "001111" => -- B7 / casella : 15
                            case sv_tipo is
                                when "0000" => B7 <= empty_L ; -- vuoto bianco
                                when "0001" => B7 <= pawn_L  ; -- pedone bianco
                                when "0010" => B7 <= king_L  ; -- re bianco
                                when "0011" => B7 <= queen_L ; -- regina bianco
                                when "0100" => B7 <= bishop_L; -- alfiere bianco
                                when "0101" => B7 <= tower_L ; -- torre bianco
                                when "0110" => B7 <= horse_L ; -- cavallo bianco
                                when "1000" => B7 <= empty_D ; -- vuoto bianco  
                                when "1001" => B7 <= pawn_D  ; -- pedone nero 
                                when "1010" => B7 <= king_D  ; -- re nero     
                                when "1011" => B7 <= queen_D ; -- regina nero 
                                when "1100" => B7 <= bishop_D; -- alfiere nero
                                when "1101" => B7 <= tower_D ; -- torre nero  
                                when "1110" => B7 <= horse_D ; -- cavallo nero
                                when others => B7 <= empty_L ; -- vuoto bianco default
                            end case;
                        when "010000" => -- C0 / casella : 16
                            case sv_tipo is
                                when "0000" => C0 <= empty_L ; -- vuoto bianco
                                when "0001" => C0 <= pawn_L  ; -- pedone bianco
                                when "0010" => C0 <= king_L  ; -- re bianco
                                when "0011" => C0 <= queen_L ; -- regina bianco
                                when "0100" => C0 <= bishop_L; -- alfiere bianco
                                when "0101" => C0 <= tower_L ; -- torre bianco
                                when "0110" => C0 <= horse_L ; -- cavallo bianco
                                when "1000" => C0 <= empty_D ; -- vuoto bianco  
                                when "1001" => C0 <= pawn_D  ; -- pedone nero 
                                when "1010" => C0 <= king_D  ; -- re nero     
                                when "1011" => C0 <= queen_D ; -- regina nero 
                                when "1100" => C0 <= bishop_D; -- alfiere nero
                                when "1101" => C0 <= tower_D ; -- torre nero  
                                when "1110" => C0 <= horse_D ; -- cavallo nero
                                when others => C0 <= empty_L ; -- vuoto bianco default
                            end case;
                        when "010001" => -- C1 / casella : 17
                            case sv_tipo is
                                when "0000" => C1 <= empty_L ; -- vuoto bianco
                                when "0001" => C1 <= pawn_L  ; -- pedone bianco
                                when "0010" => C1 <= king_L  ; -- re bianco
                                when "0011" => C1 <= queen_L ; -- regina bianco
                                when "0100" => C1 <= bishop_L; -- alfiere bianco
                                when "0101" => C1 <= tower_L ; -- torre bianco
                                when "0110" => C1 <= horse_L ; -- cavallo bianco
                                when "1000" => C1 <= empty_D ; -- vuoto bianco  
                                when "1001" => C1 <= pawn_D  ; -- pedone nero 
                                when "1010" => C1 <= king_D  ; -- re nero     
                                when "1011" => C1 <= queen_D ; -- regina nero 
                                when "1100" => C1 <= bishop_D; -- alfiere nero
                                when "1101" => C1 <= tower_D ; -- torre nero  
                                when "1110" => C1 <= horse_D ; -- cavallo nero
                                when others => C1 <= empty_L ; -- vuoto bianco default
                            end case;
                        when "010010" => -- C2 / casella : 18
                            case sv_tipo is
                                when "0000" => C2 <= empty_L ; -- vuoto bianco
                                when "0001" => C2 <= pawn_L  ; -- pedone bianco
                                when "0010" => C2 <= king_L  ; -- re bianco
                                when "0011" => C2 <= queen_L ; -- regina bianco
                                when "0100" => C2 <= bishop_L; -- alfiere bianco
                                when "0101" => C2 <= tower_L ; -- torre bianco
                                when "0110" => C2 <= horse_L ; -- cavallo bianco
                                when "1000" => C2 <= empty_D ; -- vuoto bianco  
                                when "1001" => C2 <= pawn_D  ; -- pedone nero 
                                when "1010" => C2 <= king_D  ; -- re nero     
                                when "1011" => C2 <= queen_D ; -- regina nero 
                                when "1100" => C2 <= bishop_D; -- alfiere nero
                                when "1101" => C2 <= tower_D ; -- torre nero  
                                when "1110" => C2 <= horse_D ; -- cavallo nero
                                when others => C2 <= empty_L ; -- vuoto bianco default
                            end case;
                        when "010011" => -- C3 / casella : 19
                            case sv_tipo is
                                when "0000" => C3 <= empty_L ; -- vuoto bianco
                                when "0001" => C3 <= pawn_L  ; -- pedone bianco
                                when "0010" => C3 <= king_L  ; -- re bianco
                                when "0011" => C3 <= queen_L ; -- regina bianco
                                when "0100" => C3 <= bishop_L; -- alfiere bianco
                                when "0101" => C3 <= tower_L ; -- torre bianco
                                when "0110" => C3 <= horse_L ; -- cavallo bianco
                                when "1000" => C3 <= empty_D ; -- vuoto bianco  
                                when "1001" => C3 <= pawn_D  ; -- pedone nero 
                                when "1010" => C3 <= king_D  ; -- re nero     
                                when "1011" => C3 <= queen_D ; -- regina nero 
                                when "1100" => C3 <= bishop_D; -- alfiere nero
                                when "1101" => C3 <= tower_D ; -- torre nero  
                                when "1110" => C3 <= horse_D ; -- cavallo nero
                                when others => C3 <= empty_L ; -- vuoto bianco default
                            end case;
                        when "010100" => -- C4 / casella : 20
                            case sv_tipo is
                                when "0000" => C4 <= empty_L ; -- vuoto bianco
                                when "0001" => C4 <= pawn_L  ; -- pedone bianco
                                when "0010" => C4 <= king_L  ; -- re bianco
                                when "0011" => C4 <= queen_L ; -- regina bianco
                                when "0100" => C4 <= bishop_L; -- alfiere bianco
                                when "0101" => C4 <= tower_L ; -- torre bianco
                                when "0110" => C4 <= horse_L ; -- cavallo bianco
                                when "1000" => C4 <= empty_D ; -- vuoto bianco  
                                when "1001" => C4 <= pawn_D  ; -- pedone nero 
                                when "1010" => C4 <= king_D  ; -- re nero     
                                when "1011" => C4 <= queen_D ; -- regina nero 
                                when "1100" => C4 <= bishop_D; -- alfiere nero
                                when "1101" => C4 <= tower_D ; -- torre nero  
                                when "1110" => C4 <= horse_D ; -- cavallo nero
                                when others => C4 <= empty_L ; -- vuoto bianco default
                            end case;
                        when "010101" => -- C5 / casella : 21
                            case sv_tipo is
                                when "0000" => C5 <= empty_L ; -- vuoto bianco
                                when "0001" => C5 <= pawn_L  ; -- pedone bianco
                                when "0010" => C5 <= king_L  ; -- re bianco
                                when "0011" => C5 <= queen_L ; -- regina bianco
                                when "0100" => C5 <= bishop_L; -- alfiere bianco
                                when "0101" => C5 <= tower_L ; -- torre bianco
                                when "0110" => C5 <= horse_L ; -- cavallo bianco
                                when "1000" => C5 <= empty_D ; -- vuoto bianco  
                                when "1001" => C5 <= pawn_D  ; -- pedone nero 
                                when "1010" => C5 <= king_D  ; -- re nero     
                                when "1011" => C5 <= queen_D ; -- regina nero 
                                when "1100" => C5 <= bishop_D; -- alfiere nero
                                when "1101" => C5 <= tower_D ; -- torre nero  
                                when "1110" => C5 <= horse_D ; -- cavallo nero
                                when others => C5 <= empty_L ; -- vuoto bianco default
                            end case;
                        when "010110" => -- C6 / casella : 22
                            case sv_tipo is
                                when "0000" => C6 <= empty_L ; -- vuoto bianco
                                when "0001" => C6 <= pawn_L  ; -- pedone bianco
                                when "0010" => C6 <= king_L  ; -- re bianco
                                when "0011" => C6 <= queen_L ; -- regina bianco
                                when "0100" => C6 <= bishop_L; -- alfiere bianco
                                when "0101" => C6 <= tower_L ; -- torre bianco
                                when "0110" => C6 <= horse_L ; -- cavallo bianco
                                when "1000" => C6 <= empty_D ; -- vuoto bianco  
                                when "1001" => C6 <= pawn_D  ; -- pedone nero 
                                when "1010" => C6 <= king_D  ; -- re nero     
                                when "1011" => C6 <= queen_D ; -- regina nero 
                                when "1100" => C6 <= bishop_D; -- alfiere nero
                                when "1101" => C6 <= tower_D ; -- torre nero  
                                when "1110" => C6 <= horse_D ; -- cavallo nero
                                when others => C6 <= empty_L ; -- vuoto bianco default
                            end case;
                        when "010111" => -- C7 / casella : 23
                            case sv_tipo is
                                when "0000" => C7 <= empty_L ; -- vuoto bianco
                                when "0001" => C7 <= pawn_L  ; -- pedone bianco
                                when "0010" => C7 <= king_L  ; -- re bianco
                                when "0011" => C7 <= queen_L ; -- regina bianco
                                when "0100" => C7 <= bishop_L; -- alfiere bianco
                                when "0101" => C7 <= tower_L ; -- torre bianco
                                when "0110" => C7 <= horse_L ; -- cavallo bianco
                                when "1000" => C7 <= empty_D ; -- vuoto bianco  
                                when "1001" => C7 <= pawn_D  ; -- pedone nero 
                                when "1010" => C7 <= king_D  ; -- re nero     
                                when "1011" => C7 <= queen_D ; -- regina nero 
                                when "1100" => C7 <= bishop_D; -- alfiere nero
                                when "1101" => C7 <= tower_D ; -- torre nero  
                                when "1110" => C7 <= horse_D ; -- cavallo nero
                                when others => C7 <= empty_L ; -- vuoto bianco default
                            end case;
                        when "011000" => -- D0 / casella : 24
                            case sv_tipo is
                                when "0000" => D0 <= empty_L ; -- vuoto bianco
                                when "0001" => D0 <= pawn_L  ; -- pedone bianco
                                when "0010" => D0 <= king_L  ; -- re bianco
                                when "0011" => D0 <= queen_L ; -- regina bianco
                                when "0100" => D0 <= bishop_L; -- alfiere bianco
                                when "0101" => D0 <= tower_L ; -- torre bianco
                                when "0110" => D0 <= horse_L ; -- cavallo bianco
                                when "1000" => D0 <= empty_D ; -- vuoto bianco  
                                when "1001" => D0 <= pawn_D  ; -- pedone nero 
                                when "1010" => D0 <= king_D  ; -- re nero     
                                when "1011" => D0 <= queen_D ; -- regina nero 
                                when "1100" => D0 <= bishop_D; -- alfiere nero
                                when "1101" => D0 <= tower_D ; -- torre nero  
                                when "1110" => D0 <= horse_D ; -- cavallo nero
                                when others => D0 <= empty_L ; -- vuoto bianco default
                            end case;
                        when "011001" => -- D1 / casella : 25
                            case sv_tipo is
                                when "0000" => D1 <= empty_L ; -- vuoto bianco
                                when "0001" => D1 <= pawn_L  ; -- pedone bianco
                                when "0010" => D1 <= king_L  ; -- re bianco
                                when "0011" => D1 <= queen_L ; -- regina bianco
                                when "0100" => D1 <= bishop_L; -- alfiere bianco
                                when "0101" => D1 <= tower_L ; -- torre bianco
                                when "0110" => D1 <= horse_L ; -- cavallo bianco
                                when "1000" => D1 <= empty_D ; -- vuoto bianco  
                                when "1001" => D1 <= pawn_D  ; -- pedone nero 
                                when "1010" => D1 <= king_D  ; -- re nero     
                                when "1011" => D1 <= queen_D ; -- regina nero 
                                when "1100" => D1 <= bishop_D; -- alfiere nero
                                when "1101" => D1 <= tower_D ; -- torre nero  
                                when "1110" => D1 <= horse_D ; -- cavallo nero
                                when others => D1 <= empty_L ; -- vuoto bianco default
                            end case;
                        when "011010" => -- D2 / casella : 26
                            case sv_tipo is
                                when "0000" => D2 <= empty_L ; -- vuoto bianco
                                when "0001" => D2 <= pawn_L  ; -- pedone bianco
                                when "0010" => D2 <= king_L  ; -- re bianco
                                when "0011" => D2 <= queen_L ; -- regina bianco
                                when "0100" => D2 <= bishop_L; -- alfiere bianco
                                when "0101" => D2 <= tower_L ; -- torre bianco
                                when "0110" => D2 <= horse_L ; -- cavallo bianco
                                when "1000" => D2 <= empty_D ; -- vuoto bianco  
                                when "1001" => D2 <= pawn_D  ; -- pedone nero 
                                when "1010" => D2 <= king_D  ; -- re nero     
                                when "1011" => D2 <= queen_D ; -- regina nero 
                                when "1100" => D2 <= bishop_D; -- alfiere nero
                                when "1101" => D2 <= tower_D ; -- torre nero  
                                when "1110" => D2 <= horse_D ; -- cavallo nero
                                when others => D2 <= empty_L ; -- vuoto bianco default
                            end case;
                        when "011011" => -- D3 / casella : 27
                            case sv_tipo is
                                when "0000" => D3 <= empty_L ; -- vuoto bianco
                                when "0001" => D3 <= pawn_L  ; -- pedone bianco
                                when "0010" => D3 <= king_L  ; -- re bianco
                                when "0011" => D3 <= queen_L ; -- regina bianco
                                when "0100" => D3 <= bishop_L; -- alfiere bianco
                                when "0101" => D3 <= tower_L ; -- torre bianco
                                when "0110" => D3 <= horse_L ; -- cavallo bianco
                                when "1000" => D3 <= empty_D ; -- vuoto bianco  
                                when "1001" => D3 <= pawn_D  ; -- pedone nero 
                                when "1010" => D3 <= king_D  ; -- re nero     
                                when "1011" => D3 <= queen_D ; -- regina nero 
                                when "1100" => D3 <= bishop_D; -- alfiere nero
                                when "1101" => D3 <= tower_D ; -- torre nero  
                                when "1110" => D3 <= horse_D ; -- cavallo nero
                                when others => D3 <= empty_L ; -- vuoto bianco default
                            end case;
                        when "011100" => -- D4 / casella : 28
                            case sv_tipo is
                                when "0000" => D4 <= empty_L ; -- vuoto bianco
                                when "0001" => D4 <= pawn_L  ; -- pedone bianco
                                when "0010" => D4 <= king_L  ; -- re bianco
                                when "0011" => D4 <= queen_L ; -- regina bianco
                                when "0100" => D4 <= bishop_L; -- alfiere bianco
                                when "0101" => D4 <= tower_L ; -- torre bianco
                                when "0110" => D4 <= horse_L ; -- cavallo bianco
                                when "1000" => D4 <= empty_D ; -- vuoto bianco  
                                when "1001" => D4 <= pawn_D  ; -- pedone nero 
                                when "1010" => D4 <= king_D  ; -- re nero     
                                when "1011" => D4 <= queen_D ; -- regina nero 
                                when "1100" => D4 <= bishop_D; -- alfiere nero
                                when "1101" => D4 <= tower_D ; -- torre nero  
                                when "1110" => D4 <= horse_D ; -- cavallo nero
                                when others => D4 <= empty_L ; -- vuoto bianco default
                            end case;
                        when "011101" => -- D5 / casella : 29
                            case sv_tipo is
                                when "0000" => D5 <= empty_L ; -- vuoto bianco
                                when "0001" => D5 <= pawn_L  ; -- pedone bianco
                                when "0010" => D5 <= king_L  ; -- re bianco
                                when "0011" => D5 <= queen_L ; -- regina bianco
                                when "0100" => D5 <= bishop_L; -- alfiere bianco
                                when "0101" => D5 <= tower_L ; -- torre bianco
                                when "0110" => D5 <= horse_L ; -- cavallo bianco
                                when "1000" => D5 <= empty_D ; -- vuoto bianco  
                                when "1001" => D5 <= pawn_D  ; -- pedone nero 
                                when "1010" => D5 <= king_D  ; -- re nero     
                                when "1011" => D5 <= queen_D ; -- regina nero 
                                when "1100" => D5 <= bishop_D; -- alfiere nero
                                when "1101" => D5 <= tower_D ; -- torre nero  
                                when "1110" => D5 <= horse_D ; -- cavallo nero
                                when others => D5 <= empty_L ; -- vuoto bianco default
                            end case;
                        when "011110" => -- D6 / casella : 30
                            case sv_tipo is
                                when "0000" => D6 <= empty_L ; -- vuoto bianco
                                when "0001" => D6 <= pawn_L  ; -- pedone bianco
                                when "0010" => D6 <= king_L  ; -- re bianco
                                when "0011" => D6 <= queen_L ; -- regina bianco
                                when "0100" => D6 <= bishop_L; -- alfiere bianco
                                when "0101" => D6 <= tower_L ; -- torre bianco
                                when "0110" => D6 <= horse_L ; -- cavallo bianco
                                when "1000" => D6 <= empty_D ; -- vuoto bianco  
                                when "1001" => D6 <= pawn_D  ; -- pedone nero 
                                when "1010" => D6 <= king_D  ; -- re nero     
                                when "1011" => D6 <= queen_D ; -- regina nero 
                                when "1100" => D6 <= bishop_D; -- alfiere nero
                                when "1101" => D6 <= tower_D ; -- torre nero  
                                when "1110" => D6 <= horse_D ; -- cavallo nero
                                when others => D6 <= empty_L ; -- vuoto bianco default
                            end case;
                        when "011111" => -- D7 / casella : 31
                            case sv_tipo is
                                when "0000" => D7 <= empty_L ; -- vuoto bianco
                                when "0001" => D7 <= pawn_L  ; -- pedone bianco
                                when "0010" => D7 <= king_L  ; -- re bianco
                                when "0011" => D7 <= queen_L ; -- regina bianco
                                when "0100" => D7 <= bishop_L; -- alfiere bianco
                                when "0101" => D7 <= tower_L ; -- torre bianco
                                when "0110" => D7 <= horse_L ; -- cavallo bianco
                                when "1000" => D7 <= empty_D ; -- vuoto bianco  
                                when "1001" => D7 <= pawn_D  ; -- pedone nero 
                                when "1010" => D7 <= king_D  ; -- re nero     
                                when "1011" => D7 <= queen_D ; -- regina nero 
                                when "1100" => D7 <= bishop_D; -- alfiere nero
                                when "1101" => D7 <= tower_D ; -- torre nero  
                                when "1110" => D7 <= horse_D ; -- cavallo nero
                                when others => D7 <= empty_L ; -- vuoto bianco default
                            end case;
                        when "100000" => -- E0 / casella : 32
                            case sv_tipo is
                                when "0000" => E0 <= empty_L ; -- vuoto bianco
                                when "0001" => E0 <= pawn_L  ; -- pedone bianco
                                when "0010" => E0 <= king_L  ; -- re bianco
                                when "0011" => E0 <= queen_L ; -- regina bianco
                                when "0100" => E0 <= bishop_L; -- alfiere bianco
                                when "0101" => E0 <= tower_L ; -- torre bianco
                                when "0110" => E0 <= horse_L ; -- cavallo bianco
                                when "1000" => E0 <= empty_D ; -- vuoto bianco  
                                when "1001" => E0 <= pawn_D  ; -- pedone nero 
                                when "1010" => E0 <= king_D  ; -- re nero     
                                when "1011" => E0 <= queen_D ; -- regina nero 
                                when "1100" => E0 <= bishop_D; -- alfiere nero
                                when "1101" => E0 <= tower_D ; -- torre nero  
                                when "1110" => E0 <= horse_D ; -- cavallo nero
                                when others => E0 <= empty_L ; -- vuoto bianco default
                            end case;
                        when "100001" => -- E1 / casella : 33
                            case sv_tipo is
                                when "0000" => E1 <= empty_L ; -- vuoto bianco
                                when "0001" => E1 <= pawn_L  ; -- pedone bianco
                                when "0010" => E1 <= king_L  ; -- re bianco
                                when "0011" => E1 <= queen_L ; -- regina bianco
                                when "0100" => E1 <= bishop_L; -- alfiere bianco
                                when "0101" => E1 <= tower_L ; -- torre bianco
                                when "0110" => E1 <= horse_L ; -- cavallo bianco
                                when "1000" => E1 <= empty_D ; -- vuoto bianco  
                                when "1001" => E1 <= pawn_D  ; -- pedone nero 
                                when "1010" => E1 <= king_D  ; -- re nero     
                                when "1011" => E1 <= queen_D ; -- regina nero 
                                when "1100" => E1 <= bishop_D; -- alfiere nero
                                when "1101" => E1 <= tower_D ; -- torre nero  
                                when "1110" => E1 <= horse_D ; -- cavallo nero
                                when others => E1 <= empty_L ; -- vuoto bianco default
                            end case;
                        when "100010" => -- E2 / casella : 34
                            case sv_tipo is
                                when "0000" => E2 <= empty_L ; -- vuoto bianco
                                when "0001" => E2 <= pawn_L  ; -- pedone bianco
                                when "0010" => E2 <= king_L  ; -- re bianco
                                when "0011" => E2 <= queen_L ; -- regina bianco
                                when "0100" => E2 <= bishop_L; -- alfiere bianco
                                when "0101" => E2 <= tower_L ; -- torre bianco
                                when "0110" => E2 <= horse_L ; -- cavallo bianco
                                when "1000" => E2 <= empty_D ; -- vuoto bianco  
                                when "1001" => E2 <= pawn_D  ; -- pedone nero 
                                when "1010" => E2 <= king_D  ; -- re nero     
                                when "1011" => E2 <= queen_D ; -- regina nero 
                                when "1100" => E2 <= bishop_D; -- alfiere nero
                                when "1101" => E2 <= tower_D ; -- torre nero  
                                when "1110" => E2 <= horse_D ; -- cavallo nero
                                when others => E2 <= empty_L ; -- vuoto bianco default
                            end case;
                        when "100011" => -- E3 / casella : 35
                            case sv_tipo is
                                when "0000" => E3 <= empty_L ; -- vuoto bianco
                                when "0001" => E3 <= pawn_L  ; -- pedone bianco
                                when "0010" => E3 <= king_L  ; -- re bianco
                                when "0011" => E3 <= queen_L ; -- regina bianco
                                when "0100" => E3 <= bishop_L; -- alfiere bianco
                                when "0101" => E3 <= tower_L ; -- torre bianco
                                when "0110" => E3 <= horse_L ; -- cavallo bianco
                                when "1000" => E3 <= empty_D ; -- vuoto bianco  
                                when "1001" => E3 <= pawn_D  ; -- pedone nero 
                                when "1010" => E3 <= king_D  ; -- re nero     
                                when "1011" => E3 <= queen_D ; -- regina nero 
                                when "1100" => E3 <= bishop_D; -- alfiere nero
                                when "1101" => E3 <= tower_D ; -- torre nero  
                                when "1110" => E3 <= horse_D ; -- cavallo nero
                                when others => E3 <= empty_L ; -- vuoto bianco default
                            end case;
                        when "100100" => -- E4 / casella : 36
                            case sv_tipo is
                                when "0000" => E4 <= empty_L ; -- vuoto bianco
                                when "0001" => E4 <= pawn_L  ; -- pedone bianco
                                when "0010" => E4 <= king_L  ; -- re bianco
                                when "0011" => E4 <= queen_L ; -- regina bianco
                                when "0100" => E4 <= bishop_L; -- alfiere bianco
                                when "0101" => E4 <= tower_L ; -- torre bianco
                                when "0110" => E4 <= horse_L ; -- cavallo bianco
                                when "1000" => E4 <= empty_D ; -- vuoto bianco  
                                when "1001" => E4 <= pawn_D  ; -- pedone nero 
                                when "1010" => E4 <= king_D  ; -- re nero     
                                when "1011" => E4 <= queen_D ; -- regina nero 
                                when "1100" => E4 <= bishop_D; -- alfiere nero
                                when "1101" => E4 <= tower_D ; -- torre nero  
                                when "1110" => E4 <= horse_D ; -- cavallo nero
                                when others => E4 <= empty_L ; -- vuoto bianco default
                            end case;
                        when "100101" => -- E5 / casella : 37
                            case sv_tipo is
                                when "0000" => E5 <= empty_L ; -- vuoto bianco
                                when "0001" => E5 <= pawn_L  ; -- pedone bianco
                                when "0010" => E5 <= king_L  ; -- re bianco
                                when "0011" => E5 <= queen_L ; -- regina bianco
                                when "0100" => E5 <= bishop_L; -- alfiere bianco
                                when "0101" => E5 <= tower_L ; -- torre bianco
                                when "0110" => E5 <= horse_L ; -- cavallo bianco
                                when "1000" => E5 <= empty_D ; -- vuoto bianco  
                                when "1001" => E5 <= pawn_D  ; -- pedone nero 
                                when "1010" => E5 <= king_D  ; -- re nero     
                                when "1011" => E5 <= queen_D ; -- regina nero 
                                when "1100" => E5 <= bishop_D; -- alfiere nero
                                when "1101" => E5 <= tower_D ; -- torre nero  
                                when "1110" => E5 <= horse_D ; -- cavallo nero
                                when others => E5 <= empty_L ; -- vuoto bianco default
                            end case;
                        when "100110" => -- E6 / casella : 38
                            case sv_tipo is
                                when "0000" => E6 <= empty_L ; -- vuoto bianco
                                when "0001" => E6 <= pawn_L  ; -- pedone bianco
                                when "0010" => E6 <= king_L  ; -- re bianco
                                when "0011" => E6 <= queen_L ; -- regina bianco
                                when "0100" => E6 <= bishop_L; -- alfiere bianco
                                when "0101" => E6 <= tower_L ; -- torre bianco
                                when "0110" => E6 <= horse_L ; -- cavallo bianco
                                when "1000" => E6 <= empty_D ; -- vuoto bianco  
                                when "1001" => E6 <= pawn_D  ; -- pedone nero 
                                when "1010" => E6 <= king_D  ; -- re nero     
                                when "1011" => E6 <= queen_D ; -- regina nero 
                                when "1100" => E6 <= bishop_D; -- alfiere nero
                                when "1101" => E6 <= tower_D ; -- torre nero  
                                when "1110" => E6 <= horse_D ; -- cavallo nero
                                when others => E6 <= empty_L ; -- vuoto bianco default
                            end case;
                        when "100111" => -- E7 / casella : 39
                            case sv_tipo is
                                when "0000" => E7 <= empty_L ; -- vuoto bianco
                                when "0001" => E7 <= pawn_L  ; -- pedone bianco
                                when "0010" => E7 <= king_L  ; -- re bianco
                                when "0011" => E7 <= queen_L ; -- regina bianco
                                when "0100" => E7 <= bishop_L; -- alfiere bianco
                                when "0101" => E7 <= tower_L ; -- torre bianco
                                when "0110" => E7 <= horse_L ; -- cavallo bianco
                                when "1000" => E7 <= empty_D ; -- vuoto bianco  
                                when "1001" => E7 <= pawn_D  ; -- pedone nero 
                                when "1010" => E7 <= king_D  ; -- re nero     
                                when "1011" => E7 <= queen_D ; -- regina nero 
                                when "1100" => E7 <= bishop_D; -- alfiere nero
                                when "1101" => E7 <= tower_D ; -- torre nero  
                                when "1110" => E7 <= horse_D ; -- cavallo nero
                                when others => E7 <= empty_L ; -- vuoto bianco default
                            end case;
                        when "101000" => -- F0 / casella : 40
                            case sv_tipo is
                                when "0000" => F0 <= empty_L ; -- vuoto bianco
                                when "0001" => F0 <= pawn_L  ; -- pedone bianco
                                when "0010" => F0 <= king_L  ; -- re bianco
                                when "0011" => F0 <= queen_L ; -- regina bianco
                                when "0100" => F0 <= bishop_L; -- alfiere bianco
                                when "0101" => F0 <= tower_L ; -- torre bianco
                                when "0110" => F0 <= horse_L ; -- cavallo bianco
                                when "1000" => F0 <= empty_D ; -- vuoto bianco  
                                when "1001" => F0 <= pawn_D  ; -- pedone nero 
                                when "1010" => F0 <= king_D  ; -- re nero     
                                when "1011" => F0 <= queen_D ; -- regina nero 
                                when "1100" => F0 <= bishop_D; -- alfiere nero
                                when "1101" => F0 <= tower_D ; -- torre nero  
                                when "1110" => F0 <= horse_D ; -- cavallo nero
                                when others => F0 <= empty_L ; -- vuoto bianco default
                            end case;
                        when "101001" => -- F1 / casella : 41
                            case sv_tipo is
                                when "0000" => F1 <= empty_L ; -- vuoto bianco
                                when "0001" => F1 <= pawn_L  ; -- pedone bianco
                                when "0010" => F1 <= king_L  ; -- re bianco
                                when "0011" => F1 <= queen_L ; -- regina bianco
                                when "0100" => F1 <= bishop_L; -- alfiere bianco
                                when "0101" => F1 <= tower_L ; -- torre bianco
                                when "0110" => F1 <= horse_L ; -- cavallo bianco
                                when "1000" => F1 <= empty_D ; -- vuoto bianco  
                                when "1001" => F1 <= pawn_D  ; -- pedone nero 
                                when "1010" => F1 <= king_D  ; -- re nero     
                                when "1011" => F1 <= queen_D ; -- regina nero 
                                when "1100" => F1 <= bishop_D; -- alfiere nero
                                when "1101" => F1 <= tower_D ; -- torre nero  
                                when "1110" => F1 <= horse_D ; -- cavallo nero
                                when others => F1 <= empty_L ; -- vuoto bianco default
                            end case;  
                        when "101010" => -- F2 / casella : 42
                            case sv_tipo is
                                when "0000" => F2 <= empty_L ; -- vuoto bianco
                                when "0001" => F2 <= pawn_L  ; -- pedone bianco
                                when "0010" => F2 <= king_L  ; -- re bianco
                                when "0011" => F2 <= queen_L ; -- regina bianco
                                when "0100" => F2 <= bishop_L; -- alfiere bianco
                                when "0101" => F2 <= tower_L ; -- torre bianco
                                when "0110" => F2 <= horse_L ; -- cavallo bianco
                                when "1000" => F2 <= empty_D ; -- vuoto bianco  
                                when "1001" => F2 <= pawn_D  ; -- pedone nero 
                                when "1010" => F2 <= king_D  ; -- re nero     
                                when "1011" => F2 <= queen_D ; -- regina nero 
                                when "1100" => F2 <= bishop_D; -- alfiere nero
                                when "1101" => F2 <= tower_D ; -- torre nero  
                                when "1110" => F2 <= horse_D ; -- cavallo nero
                                when others => F2 <= empty_L ; -- vuoto bianco default
                            end case;
                        when "101011" => -- F3 / casella : 43
                            case sv_tipo is
                                when "0000" => F3 <= empty_L ; -- vuoto bianco
                                when "0001" => F3 <= pawn_L  ; -- pedone bianco
                                when "0010" => F3 <= king_L  ; -- re bianco
                                when "0011" => F3 <= queen_L ; -- regina bianco
                                when "0100" => F3 <= bishop_L; -- alfiere bianco
                                when "0101" => F3 <= tower_L ; -- torre bianco
                                when "0110" => F3 <= horse_L ; -- cavallo bianco
                                when "1000" => F3 <= empty_D ; -- vuoto bianco  
                                when "1001" => F3 <= pawn_D  ; -- pedone nero 
                                when "1010" => F3 <= king_D  ; -- re nero     
                                when "1011" => F3 <= queen_D ; -- regina nero 
                                when "1100" => F3 <= bishop_D; -- alfiere nero
                                when "1101" => F3 <= tower_D ; -- torre nero  
                                when "1110" => F3 <= horse_D ; -- cavallo nero
                                when others => F3 <= empty_L ; -- vuoto bianco default
                            end case;
                        when "101100" => -- F4 / casella : 44
                            case sv_tipo is
                                when "0000" => F4 <= empty_L ; -- vuoto bianco
                                when "0001" => F4 <= pawn_L  ; -- pedone bianco
                                when "0010" => F4 <= king_L  ; -- re bianco
                                when "0011" => F4 <= queen_L ; -- regina bianco
                                when "0100" => F4 <= bishop_L; -- alfiere bianco
                                when "0101" => F4 <= tower_L ; -- torre bianco
                                when "0110" => F4 <= horse_L ; -- cavallo bianco
                                when "1000" => F4 <= empty_D ; -- vuoto bianco  
                                when "1001" => F4 <= pawn_D  ; -- pedone nero 
                                when "1010" => F4 <= king_D  ; -- re nero     
                                when "1011" => F4 <= queen_D ; -- regina nero 
                                when "1100" => F4 <= bishop_D; -- alfiere nero
                                when "1101" => F4 <= tower_D ; -- torre nero  
                                when "1110" => F4 <= horse_D ; -- cavallo nero
                                when others => F4 <= empty_L ; -- vuoto bianco default
                            end case;
                        when "101101" => -- F5 / casella : 45
                            case sv_tipo is
                                when "0000" => F5 <= empty_L ; -- vuoto bianco
                                when "0001" => F5 <= pawn_L  ; -- pedone bianco
                                when "0010" => F5 <= king_L  ; -- re bianco
                                when "0011" => F5 <= queen_L ; -- regina bianco
                                when "0100" => F5 <= bishop_L; -- alfiere bianco
                                when "0101" => F5 <= tower_L ; -- torre bianco
                                when "0110" => F5 <= horse_L ; -- cavallo bianco
                                when "1000" => F5 <= empty_D ; -- vuoto bianco  
                                when "1001" => F5 <= pawn_D  ; -- pedone nero 
                                when "1010" => F5 <= king_D  ; -- re nero     
                                when "1011" => F5 <= queen_D ; -- regina nero 
                                when "1100" => F5 <= bishop_D; -- alfiere nero
                                when "1101" => F5 <= tower_D ; -- torre nero  
                                when "1110" => F5 <= horse_D ; -- cavallo nero
                                when others => F5 <= empty_L ; -- vuoto bianco default
                            end case;
                        when "101110" => -- F6 / casella : 46
                            case sv_tipo is
                                when "0000" => F6 <= empty_L ; -- vuoto bianco
                                when "0001" => F6 <= pawn_L  ; -- pedone bianco
                                when "0010" => F6 <= king_L  ; -- re bianco
                                when "0011" => F6 <= queen_L ; -- regina bianco
                                when "0100" => F6 <= bishop_L; -- alfiere bianco
                                when "0101" => F6 <= tower_L ; -- torre bianco
                                when "0110" => F6 <= horse_L ; -- cavallo bianco
                                when "1000" => F6 <= empty_D ; -- vuoto bianco  
                                when "1001" => F6 <= pawn_D  ; -- pedone nero 
                                when "1010" => F6 <= king_D  ; -- re nero     
                                when "1011" => F6 <= queen_D ; -- regina nero 
                                when "1100" => F6 <= bishop_D; -- alfiere nero
                                when "1101" => F6 <= tower_D ; -- torre nero  
                                when "1110" => F6 <= horse_D ; -- cavallo nero
                                when others => F6 <= empty_L ; -- vuoto bianco default
                            end case;
                        when "101111" => -- F7 / casella : 47
                            case sv_tipo is
                                when "0000" => F7 <= empty_L ; -- vuoto bianco
                                when "0001" => F7 <= pawn_L  ; -- pedone bianco
                                when "0010" => F7 <= king_L  ; -- re bianco
                                when "0011" => F7 <= queen_L ; -- regina bianco
                                when "0100" => F7 <= bishop_L; -- alfiere bianco
                                when "0101" => F7 <= tower_L ; -- torre bianco
                                when "0110" => F7 <= horse_L ; -- cavallo bianco
                                when "1000" => F7 <= empty_D ; -- vuoto bianco  
                                when "1001" => F7 <= pawn_D  ; -- pedone nero 
                                when "1010" => F7 <= king_D  ; -- re nero     
                                when "1011" => F7 <= queen_D ; -- regina nero 
                                when "1100" => F7 <= bishop_D; -- alfiere nero
                                when "1101" => F7 <= tower_D ; -- torre nero  
                                when "1110" => F7 <= horse_D ; -- cavallo nero
                                when others => F7 <= empty_L ; -- vuoto bianco default
                            end case;
                        when "110000" => -- G0 / casella : 48
                            case sv_tipo is
                                when "0000" => G0 <= empty_L ; -- vuoto bianco
                                when "0001" => G0 <= pawn_L  ; -- pedone bianco
                                when "0010" => G0 <= king_L  ; -- re bianco
                                when "0011" => G0 <= queen_L ; -- regina bianco
                                when "0100" => G0 <= bishop_L; -- alfiere bianco
                                when "0101" => G0 <= tower_L ; -- torre bianco
                                when "0110" => G0 <= horse_L ; -- cavallo bianco
                                when "1000" => G0 <= empty_D ; -- vuoto bianco  
                                when "1001" => G0 <= pawn_D  ; -- pedone nero 
                                when "1010" => G0 <= king_D  ; -- re nero     
                                when "1011" => G0 <= queen_D ; -- regina nero 
                                when "1100" => G0 <= bishop_D; -- alfiere nero
                                when "1101" => G0 <= tower_D ; -- torre nero  
                                when "1110" => G0 <= horse_D ; -- cavallo nero
                                when others => G0 <= empty_L ; -- vuoto bianco default
                            end case;
                        when "110001" => -- G1 / casella : 49
                            case sv_tipo is
                                when "0000" => G1 <= empty_L ; -- vuoto bianco
                                when "0001" => G1 <= pawn_L  ; -- pedone bianco
                                when "0010" => G1 <= king_L  ; -- re bianco
                                when "0011" => G1 <= queen_L ; -- regina bianco
                                when "0100" => G1 <= bishop_L; -- alfiere bianco
                                when "0101" => G1 <= tower_L ; -- torre bianco
                                when "0110" => G1 <= horse_L ; -- cavallo bianco
                                when "1000" => G1 <= empty_D ; -- vuoto bianco  
                                when "1001" => G1 <= pawn_D  ; -- pedone nero 
                                when "1010" => G1 <= king_D  ; -- re nero     
                                when "1011" => G1 <= queen_D ; -- regina nero 
                                when "1100" => G1 <= bishop_D; -- alfiere nero
                                when "1101" => G1 <= tower_D ; -- torre nero  
                                when "1110" => G1 <= horse_D ; -- cavallo nero
                                when others => G1 <= empty_L ; -- vuoto bianco default
                            end case;
                        when "110010" => -- G2 / casella : 50
                            case sv_tipo is
                                when "0000" => G2 <= empty_L ; -- vuoto bianco
                                when "0001" => G2 <= pawn_L  ; -- pedone bianco
                                when "0010" => G2 <= king_L  ; -- re bianco
                                when "0011" => G2 <= queen_L ; -- regina bianco
                                when "0100" => G2 <= bishop_L; -- alfiere bianco
                                when "0101" => G2 <= tower_L ; -- torre bianco
                                when "0110" => G2 <= horse_L ; -- cavallo bianco
                                when "1000" => G2 <= empty_D ; -- vuoto bianco  
                                when "1001" => G2 <= pawn_D  ; -- pedone nero 
                                when "1010" => G2 <= king_D  ; -- re nero     
                                when "1011" => G2 <= queen_D ; -- regina nero 
                                when "1100" => G2 <= bishop_D; -- alfiere nero
                                when "1101" => G2 <= tower_D ; -- torre nero  
                                when "1110" => G2 <= horse_D ; -- cavallo nero
                                when others => G2 <= empty_L ; -- vuoto bianco default
                            end case;
                        when "110011" => -- G3 / casella : 51
                            case sv_tipo is
                                when "0000" => G3 <= empty_L ; -- vuoto bianco
                                when "0001" => G3 <= pawn_L  ; -- pedone bianco
                                when "0010" => G3 <= king_L  ; -- re bianco
                                when "0011" => G3 <= queen_L ; -- regina bianco
                                when "0100" => G3 <= bishop_L; -- alfiere bianco
                                when "0101" => G3 <= tower_L ; -- torre bianco
                                when "0110" => G3 <= horse_L ; -- cavallo bianco
                                when "1000" => G3 <= empty_D ; -- vuoto bianco  
                                when "1001" => G3 <= pawn_D  ; -- pedone nero 
                                when "1010" => G3 <= king_D  ; -- re nero     
                                when "1011" => G3 <= queen_D ; -- regina nero 
                                when "1100" => G3 <= bishop_D; -- alfiere nero
                                when "1101" => G3 <= tower_D ; -- torre nero  
                                when "1110" => G3 <= horse_D ; -- cavallo nero
                                when others => G3 <= empty_L ; -- vuoto bianco default
                            end case;
                        when "110100" => -- G4 / casella : 52
                            case sv_tipo is
                                when "0000" => G4 <= empty_L ; -- vuoto bianco
                                when "0001" => G4 <= pawn_L  ; -- pedone bianco
                                when "0010" => G4 <= king_L  ; -- re bianco
                                when "0011" => G4 <= queen_L ; -- regina bianco
                                when "0100" => G4 <= bishop_L; -- alfiere bianco
                                when "0101" => G4 <= tower_L ; -- torre bianco
                                when "0110" => G4 <= horse_L ; -- cavallo bianco
                                when "1000" => G4 <= empty_D ; -- vuoto bianco  
                                when "1001" => G4 <= pawn_D  ; -- pedone nero 
                                when "1010" => G4 <= king_D  ; -- re nero     
                                when "1011" => G4 <= queen_D ; -- regina nero 
                                when "1100" => G4 <= bishop_D; -- alfiere nero
                                when "1101" => G4 <= tower_D ; -- torre nero  
                                when "1110" => G4 <= horse_D ; -- cavallo nero
                                when others => G4 <= empty_L ; -- vuoto bianco default
                            end case;
                        when "110101" => -- G5 / casella : 53
                            case sv_tipo is
                                when "0000" => G5 <= empty_L ; -- vuoto bianco
                                when "0001" => G5 <= pawn_L  ; -- pedone bianco
                                when "0010" => G5 <= king_L  ; -- re bianco
                                when "0011" => G5 <= queen_L ; -- regina bianco
                                when "0100" => G5 <= bishop_L; -- alfiere bianco
                                when "0101" => G5 <= tower_L ; -- torre bianco
                                when "0110" => G5 <= horse_L ; -- cavallo bianco
                                when "1000" => G5 <= empty_D ; -- vuoto bianco  
                                when "1001" => G5 <= pawn_D  ; -- pedone nero 
                                when "1010" => G5 <= king_D  ; -- re nero     
                                when "1011" => G5 <= queen_D ; -- regina nero 
                                when "1100" => G5 <= bishop_D; -- alfiere nero
                                when "1101" => G5 <= tower_D ; -- torre nero  
                                when "1110" => G5 <= horse_D ; -- cavallo nero
                                when others => G5 <= empty_L ; -- vuoto bianco default
                            end case;
                        when "110110" => -- G6 / casella : 54
                            case sv_tipo is
                                when "0000" => G6 <= empty_L ; -- vuoto bianco
                                when "0001" => G6 <= pawn_L  ; -- pedone bianco
                                when "0010" => G6 <= king_L  ; -- re bianco
                                when "0011" => G6 <= queen_L ; -- regina bianco
                                when "0100" => G6 <= bishop_L; -- alfiere bianco
                                when "0101" => G6 <= tower_L ; -- torre bianco
                                when "0110" => G6 <= horse_L ; -- cavallo bianco
                                when "1000" => G6 <= empty_D ; -- vuoto bianco  
                                when "1001" => G6 <= pawn_D  ; -- pedone nero 
                                when "1010" => G6 <= king_D  ; -- re nero     
                                when "1011" => G6 <= queen_D ; -- regina nero 
                                when "1100" => G6 <= bishop_D; -- alfiere nero
                                when "1101" => G6 <= tower_D ; -- torre nero  
                                when "1110" => G6 <= horse_D ; -- cavallo nero
                                when others => G6 <= empty_L ; -- vuoto bianco default
                            end case;
                        when "110111" => -- G7 / casella : 55
                            case sv_tipo is
                                when "0000" => G7 <= empty_L ; -- vuoto bianco
                                when "0001" => G7 <= pawn_L  ; -- pedone bianco
                                when "0010" => G7 <= king_L  ; -- re bianco
                                when "0011" => G7 <= queen_L ; -- regina bianco
                                when "0100" => G7 <= bishop_L; -- alfiere bianco
                                when "0101" => G7 <= tower_L ; -- torre bianco
                                when "0110" => G7 <= horse_L ; -- cavallo bianco
                                when "1000" => G7 <= empty_D ; -- vuoto bianco  
                                when "1001" => G7 <= pawn_D  ; -- pedone nero 
                                when "1010" => G7 <= king_D  ; -- re nero     
                                when "1011" => G7 <= queen_D ; -- regina nero 
                                when "1100" => G7 <= bishop_D; -- alfiere nero
                                when "1101" => G7 <= tower_D ; -- torre nero  
                                when "1110" => G7 <= horse_D ; -- cavallo nero
                                when others => G7 <= empty_L ; -- vuoto bianco default
                            end case;
                        when "111000" => -- H0 / casella : 56
                            case sv_tipo is
                                when "0000" => H0 <= empty_L ; -- vuoto bianco
                                when "0001" => H0 <= pawn_L  ; -- pedone bianco
                                when "0010" => H0 <= king_L  ; -- re bianco
                                when "0011" => H0 <= queen_L ; -- regina bianco
                                when "0100" => H0 <= bishop_L; -- alfiere bianco
                                when "0101" => H0 <= tower_L ; -- torre bianco
                                when "0110" => H0 <= horse_L ; -- cavallo bianco
                                when "1000" => H0 <= empty_D ; -- vuoto bianco  
                                when "1001" => H0 <= pawn_D  ; -- pedone nero 
                                when "1010" => H0 <= king_D  ; -- re nero     
                                when "1011" => H0 <= queen_D ; -- regina nero 
                                when "1100" => H0 <= bishop_D; -- alfiere nero
                                when "1101" => H0 <= tower_D ; -- torre nero  
                                when "1110" => H0 <= horse_D ; -- cavallo nero
                                when others => H0 <= empty_L ; -- vuoto bianco default
                            end case;
                        when "111001" => -- H1 / casella : 57
                            case sv_tipo is
                                when "0000" => H1 <= empty_L ; -- vuoto bianco
                                when "0001" => H1 <= pawn_L  ; -- pedone bianco
                                when "0010" => H1 <= king_L  ; -- re bianco
                                when "0011" => H1 <= queen_L ; -- regina bianco
                                when "0100" => H1 <= bishop_L; -- alfiere bianco
                                when "0101" => H1 <= tower_L ; -- torre bianco
                                when "0110" => H1 <= horse_L ; -- cavallo bianco
                                when "1000" => H1 <= empty_D ; -- vuoto bianco  
                                when "1001" => H1 <= pawn_D  ; -- pedone nero 
                                when "1010" => H1 <= king_D  ; -- re nero     
                                when "1011" => H1 <= queen_D ; -- regina nero 
                                when "1100" => H1 <= bishop_D; -- alfiere nero
                                when "1101" => H1 <= tower_D ; -- torre nero  
                                when "1110" => H1 <= horse_D ; -- cavallo nero
                                when others => H1 <= empty_L ; -- vuoto bianco default
                            end case;
                        when "111010" => -- H2 / casella : 58
                            case sv_tipo is
                                when "0000" => H2 <= empty_L ; -- vuoto bianco
                                when "0001" => H2 <= pawn_L  ; -- pedone bianco
                                when "0010" => H2 <= king_L  ; -- re bianco
                                when "0011" => H2 <= queen_L ; -- regina bianco
                                when "0100" => H2 <= bishop_L; -- alfiere bianco
                                when "0101" => H2 <= tower_L ; -- torre bianco
                                when "0110" => H2 <= horse_L ; -- cavallo bianco
                                when "1000" => H2 <= empty_D ; -- vuoto bianco  
                                when "1001" => H2 <= pawn_D  ; -- pedone nero 
                                when "1010" => H2 <= king_D  ; -- re nero     
                                when "1011" => H2 <= queen_D ; -- regina nero 
                                when "1100" => H2 <= bishop_D; -- alfiere nero
                                when "1101" => H2 <= tower_D ; -- torre nero  
                                when "1110" => H2 <= horse_D ; -- cavallo nero
                                when others => H2 <= empty_L ; -- vuoto bianco default
                            end case;
                        when "111011" => -- H3 / casella : 59
                            case sv_tipo is
                                when "0000" => H3 <= empty_L ; -- vuoto bianco
                                when "0001" => H3 <= pawn_L  ; -- pedone bianco
                                when "0010" => H3 <= king_L  ; -- re bianco
                                when "0011" => H3 <= queen_L ; -- regina bianco
                                when "0100" => H3 <= bishop_L; -- alfiere bianco
                                when "0101" => H3 <= tower_L ; -- torre bianco
                                when "0110" => H3 <= horse_L ; -- cavallo bianco
                                when "1000" => H3 <= empty_D ; -- vuoto bianco  
                                when "1001" => H3 <= pawn_D  ; -- pedone nero 
                                when "1010" => H3 <= king_D  ; -- re nero     
                                when "1011" => H3 <= queen_D ; -- regina nero 
                                when "1100" => H3 <= bishop_D; -- alfiere nero
                                when "1101" => H3 <= tower_D ; -- torre nero  
                                when "1110" => H3 <= horse_D ; -- cavallo nero
                                when others => H3 <= empty_L ; -- vuoto bianco default
                            end case;
                        when "111100" => -- H4 / casella : 60
                            case sv_tipo is
                                when "0000" => H4 <= empty_L ; -- vuoto bianco
                                when "0001" => H4 <= pawn_L  ; -- pedone bianco
                                when "0010" => H4 <= king_L  ; -- re bianco
                                when "0011" => H4 <= queen_L ; -- regina bianco
                                when "0100" => H4 <= bishop_L; -- alfiere bianco
                                when "0101" => H4 <= tower_L ; -- torre bianco
                                when "0110" => H4 <= horse_L ; -- cavallo bianco
                                when "1000" => H4 <= empty_D ; -- vuoto bianco  
                                when "1001" => H4 <= pawn_D  ; -- pedone nero 
                                when "1010" => H4 <= king_D  ; -- re nero     
                                when "1011" => H4 <= queen_D ; -- regina nero 
                                when "1100" => H4 <= bishop_D; -- alfiere nero
                                when "1101" => H4 <= tower_D ; -- torre nero  
                                when "1110" => H4 <= horse_D ; -- cavallo nero
                                when others => H4 <= empty_L ; -- vuoto bianco default
                            end case;
                        when "111101" => -- H5 / casella : 61
                            case sv_tipo is
                                when "0000" => H5 <= empty_L ; -- vuoto bianco
                                when "0001" => H5 <= pawn_L  ; -- pedone bianco
                                when "0010" => H5 <= king_L  ; -- re bianco
                                when "0011" => H5 <= queen_L ; -- regina bianco
                                when "0100" => H5 <= bishop_L; -- alfiere bianco
                                when "0101" => H5 <= tower_L ; -- torre bianco
                                when "0110" => H5 <= horse_L ; -- cavallo bianco
                                when "1000" => H5 <= empty_D ; -- vuoto bianco  
                                when "1001" => H5 <= pawn_D  ; -- pedone nero 
                                when "1010" => H5 <= king_D  ; -- re nero     
                                when "1011" => H5 <= queen_D ; -- regina nero 
                                when "1100" => H5 <= bishop_D; -- alfiere nero
                                when "1101" => H5 <= tower_D ; -- torre nero  
                                when "1110" => H5 <= horse_D ; -- cavallo nero
                                when others => H5 <= empty_L ; -- vuoto bianco default
                            end case;
                        when "111110" => -- H6 / casella : 62
                            case sv_tipo is
                                when "0000" => H6 <= empty_L ; -- vuoto bianco
                                when "0001" => H6 <= pawn_L  ; -- pedone bianco
                                when "0010" => H6 <= king_L  ; -- re bianco
                                when "0011" => H6 <= queen_L ; -- regina bianco
                                when "0100" => H6 <= bishop_L; -- alfiere bianco
                                when "0101" => H6 <= tower_L ; -- torre bianco
                                when "0110" => H6 <= horse_L ; -- cavallo bianco
                                when "1000" => H6 <= empty_D ; -- vuoto bianco  
                                when "1001" => H6 <= pawn_D  ; -- pedone nero 
                                when "1010" => H6 <= king_D  ; -- re nero     
                                when "1011" => H6 <= queen_D ; -- regina nero 
                                when "1100" => H6 <= bishop_D; -- alfiere nero
                                when "1101" => H6 <= tower_D ; -- torre nero  
                                when "1110" => H6 <= horse_D ; -- cavallo nero
                                when others => H6 <= empty_L ; -- vuoto bianco default
                            end case;
                        when "111111" => -- H7 / casella : 63
                            case sv_tipo is
                                when "0000" => H7 <= empty_L ; -- vuoto bianco
                                when "0001" => H7 <= pawn_L  ; -- pedone bianco
                                when "0010" => H7 <= king_L  ; -- re bianco
                                when "0011" => H7 <= queen_L ; -- regina bianco
                                when "0100" => H7 <= bishop_L; -- alfiere bianco
                                when "0101" => H7 <= tower_L ; -- torre bianco
                                when "0110" => H7 <= horse_L ; -- cavallo bianco
                                when "1000" => H7 <= empty_D ; -- vuoto bianco  
                                when "1001" => H7 <= pawn_D  ; -- pedone nero 
                                when "1010" => H7 <= king_D  ; -- re nero     
                                when "1011" => H7 <= queen_D ; -- regina nero 
                                when "1100" => H7 <= bishop_D; -- alfiere nero
                                when "1101" => H7 <= tower_D ; -- torre nero  
                                when "1110" => H7 <= horse_D ; -- cavallo nero
                                when others => H7 <= empty_L ; -- vuoto bianco default
                            end case;
                        when others   => -- non ce ne sono
                            case sv_tipo is
                                when "0000" => A0 <= empty_L ; -- vuoto bianco
                                when "0001" => A0 <= pawn_L  ; -- pedone bianco
                                when "0010" => A0 <= king_L  ; -- re bianco
                                when "0011" => A0 <= queen_L ; -- regina bianco
                                when "0100" => A0 <= bishop_L; -- alfiere bianco
                                when "0101" => A0 <= tower_L ; -- torre bianco
                                when "0110" => A0 <= horse_L ; -- cavallo bianco
                                when "1000" => A0 <= empty_D ; -- vuoto bianco  
                                when "1001" => A0 <= pawn_D  ; -- pedone nero 
                                when "1010" => A0 <= king_D  ; -- re nero     
                                when "1011" => A0 <= queen_D ; -- regina nero 
                                when "1100" => A0 <= bishop_D; -- alfiere nero
                                when "1101" => A0 <= tower_D ; -- torre nero  
                                when "1110" => A0 <= horse_D ; -- cavallo nero
                                when others => A0 <= empty_L ; -- vuoto bianco default
                            end case;
                    end case;
                end if;
                end if;            
            end if;
        end process;

        AGGIORNAMENTO_COLORI:   process (FRM_i_CLK_25M) begin
            if(rising_edge(FRM_i_CLK_25M)) then
                si_curs_x <= si_curs_x_reg0;
                si_curs_y <= si_curs_y_reg0;
                    if(FRM_i_ON_STATE = '1') then
                        -- Cursore su schermo
                        st_lamp_off1    <= st_lamp_off;
                        if (((si_curs_x + si_curs_y) mod 2) = 0) then
                            st_lamp_on  <= empty_D      ;
                        else
                            st_lamp_on  <= empty_L      ;
                        end if;
                        case st_stato is
                            when IDLE =>
                                st_stato        <= LAMP_ON      ;
                            when LAMP_ON =>
                                st_cursore      <= st_lamp_on   ;
                                st_stato_dopo   <= LAMP_OFF     ;
                                st_stato        <= WAIT1        ;
                            when LAMP_OFF =>
                                st_cursore      <= st_lamp_off1 ;
                                st_stato_dopo   <= LAMP_ON      ;
                                st_stato        <= WAIT1        ;
                            when WAIT1 =>
                                ss_delay_en     <= '1'          ;
                                sv_delay_ms     <= "000111110100"; -- 500
                                st_stato        <= WAIT2        ;
                            when WAIT2 =>
                                if (ss_delay_done = '1') then
                                    st_stato    <= WAIT3        ;
                                end if;
                            when WAIT3 =>
                                ss_delay_en     <= '0'          ;
                                st_stato        <= st_stato_dopo;
                            when others =>
                                st_stato        <= IDLE         ;
                                ss_delay_en     <= '0'          ;
                        end case;
                        -- Fine cursore su schermo

                        --A0
                        if ((sv_v_cnt >= 0 and sv_v_cnt <= 19 and sv_h_cnt >= 80 and sv_h_cnt <= 139) 
                            or (sv_v_cnt >= 20 and sv_v_cnt <= 39 and sv_h_cnt >= 80 and sv_h_cnt <= 99) 
                            or (sv_v_cnt >= 20 and sv_v_cnt <= 39 and sv_h_cnt >= 120 and sv_h_cnt <= 139) 
                            or (sv_v_cnt >= 40 and sv_v_cnt <= 59 and sv_h_cnt >= 80 and sv_h_cnt <= 139)) then
                            FRM_o_R         <= "1111";
                            FRM_o_G         <= "1111";
                            FRM_o_B         <= "1111";
                        elsif (sv_v_cnt >= 20 and sv_v_cnt <= 39 and sv_h_cnt >= 100 and sv_h_cnt <= 119) then
                            sv_x_matrix     <= sv_h_cnt - 100;
                            sv_y_matrix     <= sv_v_cnt -  20;
                            if (si_curs_x = 0 and si_curs_y = 0) then
                                st_lamp_off <= A0;
                                FRM_o_R     <= st_cursore(to_integer(sv_y_matrix),to_integer(sv_x_matrix))(11 downto 8);
                                FRM_o_G     <= st_cursore(to_integer(sv_y_matrix),to_integer(sv_x_matrix))( 7 downto 4);
                                FRM_o_B     <= st_cursore(to_integer(sv_y_matrix),to_integer(sv_x_matrix))( 3 downto 0);
                            else
                                FRM_o_R     <= A0(to_integer(sv_y_matrix),to_integer(sv_x_matrix))(11 downto 8);
                                FRM_o_G     <= A0(to_integer(sv_y_matrix),to_integer(sv_x_matrix))( 7 downto 4);
                                FRM_o_B     <= A0(to_integer(sv_y_matrix),to_integer(sv_x_matrix))( 3 downto 0);
                            end if;
                            --FRM_o_R <= A0(to_integer(sv_y_matrix),to_integer(sv_x_matrix))(11 downto 8);
                            --FRM_o_G <= A0(to_integer(sv_y_matrix),to_integer(sv_x_matrix))( 7 downto 4);
                            --FRM_o_B <= A0(to_integer(sv_y_matrix),to_integer(sv_x_matrix))( 3 downto 0);
                        end if;
                        --A1
                        if ((sv_v_cnt >= 0 and sv_v_cnt <= 19 and sv_h_cnt >= 140 and sv_h_cnt <= 199) 
                            or (sv_v_cnt >= 20 and sv_v_cnt <= 39 and sv_h_cnt >= 140 and sv_h_cnt <= 159) 
                            or (sv_v_cnt >= 20 and sv_v_cnt <= 39 and sv_h_cnt >= 180 and sv_h_cnt <= 199) 
                            or (sv_v_cnt >= 40 and sv_v_cnt <= 59 and sv_h_cnt >= 140 and sv_h_cnt <= 199)) then
                            FRM_o_R         <= "0000";
                            FRM_o_G         <= "0000";
                            FRM_o_B         <= "0000";
                        elsif (sv_v_cnt >= 20 and sv_v_cnt <= 39 and sv_h_cnt >= 160 and sv_h_cnt <= 179) then
                            sv_x_matrix     <= sv_h_cnt - 160;
                            sv_y_matrix     <= sv_v_cnt -  20;
                            if (si_curs_x = 1 and si_curs_y = 0) then
                                st_lamp_off <= A1;
                                FRM_o_R     <= st_cursore(to_integer(sv_y_matrix),to_integer(sv_x_matrix))(11 downto 8);
                                FRM_o_G     <= st_cursore(to_integer(sv_y_matrix),to_integer(sv_x_matrix))( 7 downto 4);
                                FRM_o_B     <= st_cursore(to_integer(sv_y_matrix),to_integer(sv_x_matrix))( 3 downto 0);
                            else
                                FRM_o_R     <= A1(to_integer(sv_y_matrix),to_integer(sv_x_matrix))(11 downto 8);
                                FRM_o_G     <= A1(to_integer(sv_y_matrix),to_integer(sv_x_matrix))( 7 downto 4);
                                FRM_o_B     <= A1(to_integer(sv_y_matrix),to_integer(sv_x_matrix))( 3 downto 0);
                            end if;
                            --FRM_o_R <= A1(to_integer(sv_y_matrix),to_integer(sv_x_matrix))(11 downto 8);
                            --FRM_o_G <= A1(to_integer(sv_y_matrix),to_integer(sv_x_matrix))( 7 downto 4);
                            --FRM_o_B <= A1(to_integer(sv_y_matrix),to_integer(sv_x_matrix))( 3 downto 0);
                        end if;
                        --A2
                        if ((sv_v_cnt >= 0 and sv_v_cnt <= 19 and sv_h_cnt >= 200 and sv_h_cnt <= 259) 
                            or (sv_v_cnt >= 20 and sv_v_cnt <= 39 and sv_h_cnt >= 200 and sv_h_cnt <= 219) 
                            or (sv_v_cnt >= 20 and sv_v_cnt <= 39 and sv_h_cnt >= 240 and sv_h_cnt <= 259) 
                            or (sv_v_cnt >= 40 and sv_v_cnt <= 59 and sv_h_cnt >= 200 and sv_h_cnt <= 259)) then
                            FRM_o_R         <= "1111";
                            FRM_o_G         <= "1111";
                            FRM_o_B         <= "1111";
                        elsif (sv_v_cnt >= 20 and sv_v_cnt <= 39 and sv_h_cnt >= 220 and sv_h_cnt <= 239) then
                            sv_x_matrix     <= sv_h_cnt - 220;
                            sv_y_matrix     <= sv_v_cnt -  20;
                            if (si_curs_x = 2 and si_curs_y = 0) then
                                st_lamp_off <= A2;
                                FRM_o_R     <= st_cursore(to_integer(sv_y_matrix),to_integer(sv_x_matrix))(11 downto 8);
                                FRM_o_G     <= st_cursore(to_integer(sv_y_matrix),to_integer(sv_x_matrix))( 7 downto 4);
                                FRM_o_B     <= st_cursore(to_integer(sv_y_matrix),to_integer(sv_x_matrix))( 3 downto 0);
                            else
                                FRM_o_R     <= A2(to_integer(sv_y_matrix),to_integer(sv_x_matrix))(11 downto 8);
                                FRM_o_G     <= A2(to_integer(sv_y_matrix),to_integer(sv_x_matrix))( 7 downto 4);
                                FRM_o_B     <= A2(to_integer(sv_y_matrix),to_integer(sv_x_matrix))( 3 downto 0);
                            end if;
                            --FRM_o_R <= A2(to_integer(sv_y_matrix),to_integer(sv_x_matrix))(11 downto 8);
                            --FRM_o_G <= A2(to_integer(sv_y_matrix),to_integer(sv_x_matrix))( 7 downto 4);
                            --FRM_o_B <= A2(to_integer(sv_y_matrix),to_integer(sv_x_matrix))( 3 downto 0);
                        end if;
                        --A3
                        if ((sv_v_cnt >= 0 and sv_v_cnt <= 19 and sv_h_cnt >= 260 and sv_h_cnt <= 319) 
                            or (sv_v_cnt >= 20 and sv_v_cnt <= 39 and sv_h_cnt >= 260 and sv_h_cnt <= 279) 
                            or (sv_v_cnt >= 20 and sv_v_cnt <= 39 and sv_h_cnt >= 300 and sv_h_cnt <= 319) 
                            or (sv_v_cnt >= 40 and sv_v_cnt <= 59 and sv_h_cnt >= 260 and sv_h_cnt <= 319)) then
                            FRM_o_R         <= "0000";
                            FRM_o_G         <= "0000";
                            FRM_o_B         <= "0000";
                        elsif (sv_v_cnt >= 20 and sv_v_cnt <= 39 and sv_h_cnt >= 280 and sv_h_cnt <= 299) then
                            sv_x_matrix     <= sv_h_cnt - 280;
                            sv_y_matrix     <= sv_v_cnt -  20;
                            if (si_curs_x = 3 and si_curs_y = 0) then
                                st_lamp_off <= A3;
                                FRM_o_R     <= st_cursore(to_integer(sv_y_matrix),to_integer(sv_x_matrix))(11 downto 8);
                                FRM_o_G     <= st_cursore(to_integer(sv_y_matrix),to_integer(sv_x_matrix))( 7 downto 4);
                                FRM_o_B     <= st_cursore(to_integer(sv_y_matrix),to_integer(sv_x_matrix))( 3 downto 0);
                            else
                                FRM_o_R     <= A3(to_integer(sv_y_matrix),to_integer(sv_x_matrix))(11 downto 8);
                                FRM_o_G     <= A3(to_integer(sv_y_matrix),to_integer(sv_x_matrix))( 7 downto 4);
                                FRM_o_B     <= A3(to_integer(sv_y_matrix),to_integer(sv_x_matrix))( 3 downto 0);
                            end if;
                            --FRM_o_R <= A3(to_integer(sv_y_matrix),to_integer(sv_x_matrix))(11 downto 8);
                            --FRM_o_G <= A3(to_integer(sv_y_matrix),to_integer(sv_x_matrix))( 7 downto 4);
                            --FRM_o_B <= A3(to_integer(sv_y_matrix),to_integer(sv_x_matrix))( 3 downto 0);
                        end if;
                        --A4
                        if ((sv_v_cnt >= 0 and sv_v_cnt <= 19 and sv_h_cnt >= 320 and sv_h_cnt <= 379) 
                            or (sv_v_cnt >= 20 and sv_v_cnt <= 39 and sv_h_cnt >= 320 and sv_h_cnt <= 339) 
                            or (sv_v_cnt >= 20 and sv_v_cnt <= 39 and sv_h_cnt >= 360 and sv_h_cnt <= 379) 
                            or (sv_v_cnt >= 40 and sv_v_cnt <= 59 and sv_h_cnt >= 320 and sv_h_cnt <= 379)) then
                            FRM_o_R         <= "1111";
                            FRM_o_G         <= "1111";
                            FRM_o_B         <= "1111";
                        elsif (sv_v_cnt >= 20 and sv_v_cnt <= 39 and sv_h_cnt >= 340 and sv_h_cnt <= 359) then
                            sv_x_matrix     <= sv_h_cnt - 340;
                            sv_y_matrix     <= sv_v_cnt -  20;
                            if (si_curs_x = 4 and si_curs_y = 0) then
                                st_lamp_off <= A4;
                                FRM_o_R     <= st_cursore(to_integer(sv_y_matrix),to_integer(sv_x_matrix))(11 downto 8);
                                FRM_o_G     <= st_cursore(to_integer(sv_y_matrix),to_integer(sv_x_matrix))( 7 downto 4);
                                FRM_o_B     <= st_cursore(to_integer(sv_y_matrix),to_integer(sv_x_matrix))( 3 downto 0);
                            else
                                FRM_o_R     <= A4(to_integer(sv_y_matrix),to_integer(sv_x_matrix))(11 downto 8);
                                FRM_o_G     <= A4(to_integer(sv_y_matrix),to_integer(sv_x_matrix))( 7 downto 4);
                                FRM_o_B     <= A4(to_integer(sv_y_matrix),to_integer(sv_x_matrix))( 3 downto 0);
                            end if;
                            --FRM_o_R <= A4(to_integer(sv_y_matrix),to_integer(sv_x_matrix))(11 downto 8);
                            --FRM_o_G <= A4(to_integer(sv_y_matrix),to_integer(sv_x_matrix))( 7 downto 4);
                            --FRM_o_B <= A4(to_integer(sv_y_matrix),to_integer(sv_x_matrix))( 3 downto 0);
                        end if;
                        --A5
                        if ((sv_v_cnt >= 0 and sv_v_cnt <= 19 and sv_h_cnt >= 380 and sv_h_cnt <= 439) 
                            or (sv_v_cnt >= 20 and sv_v_cnt <= 39 and sv_h_cnt >= 380 and sv_h_cnt <= 399) 
                            or (sv_v_cnt >= 20 and sv_v_cnt <= 39 and sv_h_cnt >= 420 and sv_h_cnt <= 439) 
                            or (sv_v_cnt >= 40 and sv_v_cnt <= 59 and sv_h_cnt >= 380 and sv_h_cnt <= 439)) then
                            FRM_o_R         <= "0000";
                            FRM_o_G         <= "0000";
                            FRM_o_B         <= "0000";
                        elsif (sv_v_cnt >= 20 and sv_v_cnt <= 39 and sv_h_cnt >= 400 and sv_h_cnt <= 419) then
                            sv_x_matrix     <= sv_h_cnt - 400;
                            sv_y_matrix     <= sv_v_cnt -  20;
                            if (si_curs_x = 5 and si_curs_y = 0) then
                                st_lamp_off <= A5;
                                FRM_o_R     <= st_cursore(to_integer(sv_y_matrix),to_integer(sv_x_matrix))(11 downto 8);
                                FRM_o_G     <= st_cursore(to_integer(sv_y_matrix),to_integer(sv_x_matrix))( 7 downto 4);
                                FRM_o_B     <= st_cursore(to_integer(sv_y_matrix),to_integer(sv_x_matrix))( 3 downto 0);
                            else
                                FRM_o_R     <= A5(to_integer(sv_y_matrix),to_integer(sv_x_matrix))(11 downto 8);
                                FRM_o_G     <= A5(to_integer(sv_y_matrix),to_integer(sv_x_matrix))( 7 downto 4);
                                FRM_o_B     <= A5(to_integer(sv_y_matrix),to_integer(sv_x_matrix))( 3 downto 0);
                            end if;
                            --FRM_o_R <= A5(to_integer(sv_y_matrix),to_integer(sv_x_matrix))(11 downto 8);
                            --FRM_o_G <= A5(to_integer(sv_y_matrix),to_integer(sv_x_matrix))( 7 downto 4);
                            --FRM_o_B <= A5(to_integer(sv_y_matrix),to_integer(sv_x_matrix))( 3 downto 0);
                        end if;
                        --A6
                        if ((sv_v_cnt >= 0 and sv_v_cnt <= 19 and sv_h_cnt >= 440 and sv_h_cnt <= 499) 
                            or (sv_v_cnt >= 20 and sv_v_cnt <= 39 and sv_h_cnt >= 440 and sv_h_cnt <= 459) 
                            or (sv_v_cnt >= 20 and sv_v_cnt <= 39 and sv_h_cnt >= 480 and sv_h_cnt <= 499) 
                            or (sv_v_cnt >= 40 and sv_v_cnt <= 59 and sv_h_cnt >= 440 and sv_h_cnt <= 499)) then                            
                            FRM_o_R         <= "1111";
                            FRM_o_G         <= "1111";
                            FRM_o_B         <= "1111";
                        elsif (sv_v_cnt >= 20 and sv_v_cnt <= 39 and sv_h_cnt >= 460 and sv_h_cnt <= 479) then
                            sv_x_matrix     <= sv_h_cnt - 460;
                            sv_y_matrix     <= sv_v_cnt -  20;
                            if (si_curs_x = 6 and si_curs_y = 0) then
                                st_lamp_off <= A6;
                                FRM_o_R     <= st_cursore(to_integer(sv_y_matrix),to_integer(sv_x_matrix))(11 downto 8);
                                FRM_o_G     <= st_cursore(to_integer(sv_y_matrix),to_integer(sv_x_matrix))( 7 downto 4);
                                FRM_o_B     <= st_cursore(to_integer(sv_y_matrix),to_integer(sv_x_matrix))( 3 downto 0);
                            else
                                FRM_o_R     <= A6(to_integer(sv_y_matrix),to_integer(sv_x_matrix))(11 downto 8);
                                FRM_o_G     <= A6(to_integer(sv_y_matrix),to_integer(sv_x_matrix))( 7 downto 4);
                                FRM_o_B     <= A6(to_integer(sv_y_matrix),to_integer(sv_x_matrix))( 3 downto 0);
                            end if;
                            --FRM_o_R <= A6(to_integer(sv_y_matrix),to_integer(sv_x_matrix))(11 downto 8);
                            --FRM_o_G <= A6(to_integer(sv_y_matrix),to_integer(sv_x_matrix))( 7 downto 4);
                            --FRM_o_B <= A6(to_integer(sv_y_matrix),to_integer(sv_x_matrix))( 3 downto 0);
                        end if;
                        --A7
                        if ((sv_v_cnt >= 0 and sv_v_cnt <= 19 and sv_h_cnt >= 500 and sv_h_cnt <= 559) 
                            or (sv_v_cnt >= 20 and sv_v_cnt <= 39 and sv_h_cnt >= 500 and sv_h_cnt <= 519) 
                            or (sv_v_cnt >= 20 and sv_v_cnt <= 39 and sv_h_cnt >= 540 and sv_h_cnt <= 559) 
                            or (sv_v_cnt >= 40 and sv_v_cnt <= 59 and sv_h_cnt >= 500 and sv_h_cnt <= 559)) then                           
                            FRM_o_R         <= "0000";
                            FRM_o_G         <= "0000";
                            FRM_o_B         <= "0000";
                        elsif (sv_v_cnt >= 20 and sv_v_cnt <= 39 and sv_h_cnt >= 520 and sv_h_cnt <= 539) then
                            sv_x_matrix     <= sv_h_cnt - 520;
                            sv_y_matrix     <= sv_v_cnt -  20;
                            if (si_curs_x = 7 and si_curs_y = 0) then
                                st_lamp_off <= A7;
                                FRM_o_R     <= st_cursore(to_integer(sv_y_matrix),to_integer(sv_x_matrix))(11 downto 8);
                                FRM_o_G     <= st_cursore(to_integer(sv_y_matrix),to_integer(sv_x_matrix))( 7 downto 4);
                                FRM_o_B     <= st_cursore(to_integer(sv_y_matrix),to_integer(sv_x_matrix))( 3 downto 0);
                            else
                                FRM_o_R     <= A7(to_integer(sv_y_matrix),to_integer(sv_x_matrix))(11 downto 8);
                                FRM_o_G     <= A7(to_integer(sv_y_matrix),to_integer(sv_x_matrix))( 7 downto 4);
                                FRM_o_B     <= A7(to_integer(sv_y_matrix),to_integer(sv_x_matrix))( 3 downto 0);
                            end if;
                            --FRM_o_R <= A7(to_integer(sv_y_matrix),to_integer(sv_x_matrix))(11 downto 8);
                            --FRM_o_G <= A7(to_integer(sv_y_matrix),to_integer(sv_x_matrix))( 7 downto 4);
                            --FRM_o_B <= A7(to_integer(sv_y_matrix),to_integer(sv_x_matrix))( 3 downto 0);
                        end if;
                        --B0
                        if ((sv_v_cnt >= 60 and sv_v_cnt <= 79 and sv_h_cnt >= 80 and sv_h_cnt <= 139) 
                            or (sv_v_cnt >= 80 and sv_v_cnt <= 99 and sv_h_cnt >= 80 and sv_h_cnt <= 99) 
                            or (sv_v_cnt >= 80 and sv_v_cnt <= 99 and sv_h_cnt >= 120 and sv_h_cnt <= 139) 
                            or (sv_v_cnt >= 100 and sv_v_cnt <= 119 and sv_h_cnt >= 80 and sv_h_cnt <= 139)) then
                            FRM_o_R         <= "0000";
                            FRM_o_G         <= "0000";
                            FRM_o_B         <= "0000";
                        elsif (sv_v_cnt >= 80 and sv_v_cnt <= 99 and sv_h_cnt >= 100 and sv_h_cnt <= 119) then
                            sv_x_matrix     <= sv_h_cnt - 100;
                            sv_y_matrix     <= sv_v_cnt -  80;
                            if (si_curs_x = 0 and si_curs_y = 1) then
                                st_lamp_off <= B0;
                                FRM_o_R     <= st_cursore(to_integer(sv_y_matrix),to_integer(sv_x_matrix))(11 downto 8);
                                FRM_o_G     <= st_cursore(to_integer(sv_y_matrix),to_integer(sv_x_matrix))( 7 downto 4);
                                FRM_o_B     <= st_cursore(to_integer(sv_y_matrix),to_integer(sv_x_matrix))( 3 downto 0);
                            else
                                FRM_o_R     <= B0(to_integer(sv_y_matrix),to_integer(sv_x_matrix))(11 downto 8);
                                FRM_o_G     <= B0(to_integer(sv_y_matrix),to_integer(sv_x_matrix))( 7 downto 4);
                                FRM_o_B     <= B0(to_integer(sv_y_matrix),to_integer(sv_x_matrix))( 3 downto 0);
                            end if;
                            --FRM_o_R <= B0(to_integer(sv_y_matrix),to_integer(sv_x_matrix))(11 downto 8);
                            --FRM_o_G <= B0(to_integer(sv_y_matrix),to_integer(sv_x_matrix))( 7 downto 4);
                            --FRM_o_B <= B0(to_integer(sv_y_matrix),to_integer(sv_x_matrix))( 3 downto 0);
                        end if;
                        --B1
                        if ((sv_v_cnt >= 60 and sv_v_cnt <= 79 and sv_h_cnt >= 140 and sv_h_cnt <= 199) 
                            or (sv_v_cnt >= 80 and sv_v_cnt <= 99 and sv_h_cnt >= 140 and sv_h_cnt <= 159) 
                            or (sv_v_cnt >= 80 and sv_v_cnt <= 99 and sv_h_cnt >= 180 and sv_h_cnt <= 199) 
                            or (sv_v_cnt >= 100 and sv_v_cnt <= 119 and sv_h_cnt >= 140 and sv_h_cnt <= 199)) then                            
                            FRM_o_R         <= "1111";
                            FRM_o_G         <= "1111";
                            FRM_o_B         <= "1111";
                        elsif (sv_v_cnt >= 80 and sv_v_cnt <= 99 and sv_h_cnt >= 160 and sv_h_cnt <= 179) then
                            sv_x_matrix     <= sv_h_cnt - 160;
                            sv_y_matrix     <= sv_v_cnt -  80;
                            if (si_curs_x = 1 and si_curs_y = 1) then
                                st_lamp_off <= B1;
                                FRM_o_R     <= st_cursore(to_integer(sv_y_matrix),to_integer(sv_x_matrix))(11 downto 8);
                                FRM_o_G     <= st_cursore(to_integer(sv_y_matrix),to_integer(sv_x_matrix))( 7 downto 4);
                                FRM_o_B     <= st_cursore(to_integer(sv_y_matrix),to_integer(sv_x_matrix))( 3 downto 0);
                            else
                                FRM_o_R     <= B1(to_integer(sv_y_matrix),to_integer(sv_x_matrix))(11 downto 8);
                                FRM_o_G     <= B1(to_integer(sv_y_matrix),to_integer(sv_x_matrix))( 7 downto 4);
                                FRM_o_B     <= B1(to_integer(sv_y_matrix),to_integer(sv_x_matrix))( 3 downto 0);
                            end if;
                            --FRM_o_R         <= B1(to_integer(sv_y_matrix),to_integer(sv_x_matrix))(11 downto 8);
                            --FRM_o_G         <= B1(to_integer(sv_y_matrix),to_integer(sv_x_matrix))( 7 downto 4);
                            --FRM_o_B         <= B1(to_integer(sv_y_matrix),to_integer(sv_x_matrix))( 3 downto 0);
                        end if;
                        --B2
                        if ((sv_v_cnt >= 60 and sv_v_cnt <= 79 and sv_h_cnt >= 200 and sv_h_cnt <= 259) 
                            or (sv_v_cnt >= 80 and sv_v_cnt <= 99 and sv_h_cnt >= 200 and sv_h_cnt <= 219) 
                            or (sv_v_cnt >= 80 and sv_v_cnt <= 99 and sv_h_cnt >= 240 and sv_h_cnt <= 259) 
                            or (sv_v_cnt >= 100 and sv_v_cnt <= 119 and sv_h_cnt >= 200 and sv_h_cnt <= 259)) then
                            FRM_o_R         <= "0000";
                            FRM_o_G         <= "0000";
                            FRM_o_B         <= "0000";
                        elsif (sv_v_cnt >= 80 and sv_v_cnt <= 99 and sv_h_cnt >= 220 and sv_h_cnt <= 239) then
                            sv_x_matrix <= sv_h_cnt - 220;
                            sv_y_matrix <= sv_v_cnt -  80;
                            if (si_curs_x = 2 and si_curs_y = 1) then
                                st_lamp_off <= B2;
                                FRM_o_R     <= st_cursore(to_integer(sv_y_matrix),to_integer(sv_x_matrix))(11 downto 8);
                                FRM_o_G     <= st_cursore(to_integer(sv_y_matrix),to_integer(sv_x_matrix))( 7 downto 4);
                                FRM_o_B     <= st_cursore(to_integer(sv_y_matrix),to_integer(sv_x_matrix))( 3 downto 0);
                            else
                                FRM_o_R     <= B2(to_integer(sv_y_matrix),to_integer(sv_x_matrix))(11 downto 8);
                                FRM_o_G     <= B2(to_integer(sv_y_matrix),to_integer(sv_x_matrix))( 7 downto 4);
                                FRM_o_B     <= B2(to_integer(sv_y_matrix),to_integer(sv_x_matrix))( 3 downto 0);
                            end if;
                            --FRM_o_R <= B2(to_integer(sv_y_matrix),to_integer(sv_x_matrix))(11 downto 8);
                            --FRM_o_G <= B2(to_integer(sv_y_matrix),to_integer(sv_x_matrix))( 7 downto 4);
                            --FRM_o_B <= B2(to_integer(sv_y_matrix),to_integer(sv_x_matrix))( 3 downto 0);
                        end if;
                        --B3
                        if ((sv_v_cnt >= 60 and sv_v_cnt <= 79 and sv_h_cnt >= 260 and sv_h_cnt <= 319) 
                            or (sv_v_cnt >= 80 and sv_v_cnt <= 99 and sv_h_cnt >= 260 and sv_h_cnt <= 279) 
                            or (sv_v_cnt >= 80 and sv_v_cnt <= 99 and sv_h_cnt >= 300 and sv_h_cnt <= 319) 
                            or (sv_v_cnt >= 100 and sv_v_cnt <= 119 and sv_h_cnt >= 260 and sv_h_cnt <= 319)) then
                            FRM_o_R <= "1111";
                            FRM_o_G <= "1111";
                            FRM_o_B <= "1111";
                        elsif (sv_v_cnt >= 80 and sv_v_cnt <= 99 and sv_h_cnt >= 280 and sv_h_cnt <= 299) then
                            sv_x_matrix <= sv_h_cnt - 280;
                            sv_y_matrix <= sv_v_cnt -  80;
                            if (si_curs_x = 3 and si_curs_y = 1) then
                                st_lamp_off <= B3;
                                FRM_o_R     <= st_cursore(to_integer(sv_y_matrix),to_integer(sv_x_matrix))(11 downto 8);
                                FRM_o_G     <= st_cursore(to_integer(sv_y_matrix),to_integer(sv_x_matrix))( 7 downto 4);
                                FRM_o_B     <= st_cursore(to_integer(sv_y_matrix),to_integer(sv_x_matrix))( 3 downto 0);
                            else
                                FRM_o_R     <= B3(to_integer(sv_y_matrix),to_integer(sv_x_matrix))(11 downto 8);
                                FRM_o_G     <= B3(to_integer(sv_y_matrix),to_integer(sv_x_matrix))( 7 downto 4);
                                FRM_o_B     <= B3(to_integer(sv_y_matrix),to_integer(sv_x_matrix))( 3 downto 0);
                            end if;
                            --FRM_o_R <= B3(to_integer(sv_y_matrix),to_integer(sv_x_matrix))(11 downto 8);
                            --FRM_o_G <= B3(to_integer(sv_y_matrix),to_integer(sv_x_matrix))( 7 downto 4);
                            --FRM_o_B <= B3(to_integer(sv_y_matrix),to_integer(sv_x_matrix))( 3 downto 0);
                        end if;
                        --B4
                        if ((sv_v_cnt >= 60 and sv_v_cnt <= 79 and sv_h_cnt >= 320 and sv_h_cnt <= 379) 
                            or (sv_v_cnt >= 80 and sv_v_cnt <= 99 and sv_h_cnt >= 320 and sv_h_cnt <= 339) 
                            or (sv_v_cnt >= 80 and sv_v_cnt <= 99 and sv_h_cnt >= 360 and sv_h_cnt <= 379) 
                            or (sv_v_cnt >= 100 and sv_v_cnt <= 119 and sv_h_cnt >= 320 and sv_h_cnt <= 379)) then
                            FRM_o_R <= "0000";
                            FRM_o_G <= "0000";
                            FRM_o_B <= "0000";
                        elsif (sv_v_cnt >= 80 and sv_v_cnt <= 99 and sv_h_cnt >= 340 and sv_h_cnt <= 359) then
                            sv_x_matrix <= sv_h_cnt - 340;
                            sv_y_matrix <= sv_v_cnt -  80;
                            if (si_curs_x = 4 and si_curs_y = 1) then
                                st_lamp_off <= B4;
                                FRM_o_R     <= st_cursore(to_integer(sv_y_matrix),to_integer(sv_x_matrix))(11 downto 8);
                                FRM_o_G     <= st_cursore(to_integer(sv_y_matrix),to_integer(sv_x_matrix))( 7 downto 4);
                                FRM_o_B     <= st_cursore(to_integer(sv_y_matrix),to_integer(sv_x_matrix))( 3 downto 0);
                            else
                                FRM_o_R     <= B4(to_integer(sv_y_matrix),to_integer(sv_x_matrix))(11 downto 8);
                                FRM_o_G     <= B4(to_integer(sv_y_matrix),to_integer(sv_x_matrix))( 7 downto 4);
                                FRM_o_B     <= B4(to_integer(sv_y_matrix),to_integer(sv_x_matrix))( 3 downto 0);
                            end if;
                            --FRM_o_R <= B4(to_integer(sv_y_matrix),to_integer(sv_x_matrix))(11 downto 8);
                            --FRM_o_G <= B4(to_integer(sv_y_matrix),to_integer(sv_x_matrix))( 7 downto 4);
                            --FRM_o_B <= B4(to_integer(sv_y_matrix),to_integer(sv_x_matrix))( 3 downto 0);+
                        end if;
                        --B5
                        if ((sv_v_cnt >= 60 and sv_v_cnt <= 79 and sv_h_cnt >= 380 and sv_h_cnt <= 439) 
                            or (sv_v_cnt >= 80 and sv_v_cnt <= 99 and sv_h_cnt >= 380 and sv_h_cnt <= 399) 
                            or (sv_v_cnt >= 80 and sv_v_cnt <= 99 and sv_h_cnt >= 420 and sv_h_cnt <= 439) 
                            or (sv_v_cnt >= 100 and sv_v_cnt <= 119 and sv_h_cnt >= 380 and sv_h_cnt <= 439)) then
                            FRM_o_R <= "1111";
                            FRM_o_G <= "1111";
                            FRM_o_B <= "1111";
                        elsif (sv_v_cnt >= 80 and sv_v_cnt <= 99 and sv_h_cnt >= 400 and sv_h_cnt <= 419) then
                            sv_x_matrix <= sv_h_cnt - 400;
                            sv_y_matrix <= sv_v_cnt -  80;
                            if (si_curs_x = 5 and si_curs_y = 1) then
                                st_lamp_off <= B5;
                                FRM_o_R     <= st_cursore(to_integer(sv_y_matrix),to_integer(sv_x_matrix))(11 downto 8);
                                FRM_o_G     <= st_cursore(to_integer(sv_y_matrix),to_integer(sv_x_matrix))( 7 downto 4);
                                FRM_o_B     <= st_cursore(to_integer(sv_y_matrix),to_integer(sv_x_matrix))( 3 downto 0);
                            else
                                FRM_o_R     <= B5(to_integer(sv_y_matrix),to_integer(sv_x_matrix))(11 downto 8);
                                FRM_o_G     <= B5(to_integer(sv_y_matrix),to_integer(sv_x_matrix))( 7 downto 4);
                                FRM_o_B     <= B5(to_integer(sv_y_matrix),to_integer(sv_x_matrix))( 3 downto 0);
                            end if;
                            --FRM_o_R <= B5(to_integer(sv_y_matrix),to_integer(sv_x_matrix))(11 downto 8);
                            --FRM_o_G <= B5(to_integer(sv_y_matrix),to_integer(sv_x_matrix))( 7 downto 4);
                            --FRM_o_B <= B5(to_integer(sv_y_matrix),to_integer(sv_x_matrix))( 3 downto 0);
                        end if;
                        --B6
                        if ((sv_v_cnt >= 60 and sv_v_cnt <= 79 and sv_h_cnt >= 440 and sv_h_cnt <= 499) 
                            or (sv_v_cnt >= 80 and sv_v_cnt <= 99 and sv_h_cnt >= 440 and sv_h_cnt <= 459) 
                            or (sv_v_cnt >= 80 and sv_v_cnt <= 99 and sv_h_cnt >= 480 and sv_h_cnt <= 499) 
                            or (sv_v_cnt >= 100 and sv_v_cnt <= 119 and sv_h_cnt >= 440 and sv_h_cnt <= 499)) then
                            FRM_o_R <= "0000";
                            FRM_o_G <= "0000";
                            FRM_o_B <= "0000";
                        elsif (sv_v_cnt >= 80 and sv_v_cnt <= 99 and sv_h_cnt >= 460 and sv_h_cnt <= 479) then
                            sv_x_matrix <= sv_h_cnt - 460;
                            sv_y_matrix <= sv_v_cnt -  80;
                            if (si_curs_x = 6 and si_curs_y = 1) then
                                st_lamp_off <= B6;
                                FRM_o_R     <= st_cursore(to_integer(sv_y_matrix),to_integer(sv_x_matrix))(11 downto 8);
                                FRM_o_G     <= st_cursore(to_integer(sv_y_matrix),to_integer(sv_x_matrix))( 7 downto 4);
                                FRM_o_B     <= st_cursore(to_integer(sv_y_matrix),to_integer(sv_x_matrix))( 3 downto 0);
                            else
                                FRM_o_R     <= B6(to_integer(sv_y_matrix),to_integer(sv_x_matrix))(11 downto 8);
                                FRM_o_G     <= B6(to_integer(sv_y_matrix),to_integer(sv_x_matrix))( 7 downto 4);
                                FRM_o_B     <= B6(to_integer(sv_y_matrix),to_integer(sv_x_matrix))( 3 downto 0);
                            end if;
                            --FRM_o_R <= B6(to_integer(sv_y_matrix),to_integer(sv_x_matrix))(11 downto 8);
                            --FRM_o_G <= B6(to_integer(sv_y_matrix),to_integer(sv_x_matrix))( 7 downto 4);
                            --FRM_o_B <= B6(to_integer(sv_y_matrix),to_integer(sv_x_matrix))( 3 downto 0);
                        end if;
                        --B7
                        if ((sv_v_cnt >= 60 and sv_v_cnt <= 79 and sv_h_cnt >= 500 and sv_h_cnt <= 559) 
                            or (sv_v_cnt >= 80 and sv_v_cnt <= 99 and sv_h_cnt >= 500 and sv_h_cnt <= 519) 
                            or (sv_v_cnt >= 80 and sv_v_cnt <= 99 and sv_h_cnt >= 540 and sv_h_cnt <= 559) 
                            or (sv_v_cnt >= 100 and sv_v_cnt <= 119 and sv_h_cnt >= 500 and sv_h_cnt <= 559)) then
                            FRM_o_R <= "1111";
                            FRM_o_G <= "1111";
                            FRM_o_B <= "1111";
                        elsif (sv_v_cnt >= 80 and sv_v_cnt <= 119 and sv_h_cnt >= 520 and sv_h_cnt <= 539) then
                            sv_x_matrix <= sv_h_cnt - 520;
                            sv_y_matrix <= sv_v_cnt -  80;
                            if (si_curs_x = 7 and si_curs_y = 1) then
                                st_lamp_off <= B7;
                                FRM_o_R     <= st_cursore(to_integer(sv_y_matrix),to_integer(sv_x_matrix))(11 downto 8);
                                FRM_o_G     <= st_cursore(to_integer(sv_y_matrix),to_integer(sv_x_matrix))( 7 downto 4);
                                FRM_o_B     <= st_cursore(to_integer(sv_y_matrix),to_integer(sv_x_matrix))( 3 downto 0);
                            else
                                FRM_o_R     <= B7(to_integer(sv_y_matrix),to_integer(sv_x_matrix))(11 downto 8);
                                FRM_o_G     <= B7(to_integer(sv_y_matrix),to_integer(sv_x_matrix))( 7 downto 4);
                                FRM_o_B     <= B7(to_integer(sv_y_matrix),to_integer(sv_x_matrix))( 3 downto 0);
                            end if;
                            --FRM_o_R <= B7(to_integer(sv_y_matrix),to_integer(sv_x_matrix))(11 downto 8);
                            --FRM_o_G <= B7(to_integer(sv_y_matrix),to_integer(sv_x_matrix))( 7 downto 4);
                            --FRM_o_B <= B7(to_integer(sv_y_matrix),to_integer(sv_x_matrix))( 3 downto 0);
                        end if;
                        --C0
                        if ((sv_v_cnt >= 120 and sv_v_cnt <= 139 and sv_h_cnt >= 80 and sv_h_cnt <= 139) 
                            or (sv_v_cnt >= 140 and sv_v_cnt <= 159 and sv_h_cnt >= 80 and sv_h_cnt <= 99) 
                            or (sv_v_cnt >= 140 and sv_v_cnt <= 159 and sv_h_cnt >= 120 and sv_h_cnt <= 139) 
                            or (sv_v_cnt >= 160 and sv_v_cnt <= 179 and sv_h_cnt >= 80 and sv_h_cnt <= 139)) then
                            FRM_o_R <= "1111";
                            FRM_o_G <= "1111";
                            FRM_o_B <= "1111";
                        elsif (sv_v_cnt >= 140 and sv_v_cnt <= 159 and sv_h_cnt >= 100 and sv_h_cnt <= 119) then
                            sv_x_matrix <= sv_h_cnt - 100;
                            sv_y_matrix <= sv_v_cnt - 140;
                            if (si_curs_x = 0 and si_curs_y = 2) then
                                st_lamp_off <= C0;
                                FRM_o_R     <= st_cursore(to_integer(sv_y_matrix),to_integer(sv_x_matrix))(11 downto 8);
                                FRM_o_G     <= st_cursore(to_integer(sv_y_matrix),to_integer(sv_x_matrix))( 7 downto 4);
                                FRM_o_B     <= st_cursore(to_integer(sv_y_matrix),to_integer(sv_x_matrix))( 3 downto 0);
                            else
                                FRM_o_R     <= C0(to_integer(sv_y_matrix),to_integer(sv_x_matrix))(11 downto 8);
                                FRM_o_G     <= C0(to_integer(sv_y_matrix),to_integer(sv_x_matrix))( 7 downto 4);
                                FRM_o_B     <= C0(to_integer(sv_y_matrix),to_integer(sv_x_matrix))( 3 downto 0);
                            end if;
                            --FRM_o_R <= C0(to_integer(sv_y_matrix),to_integer(sv_x_matrix))(11 downto 8);
                            --FRM_o_G <= C0(to_integer(sv_y_matrix),to_integer(sv_x_matrix))( 7 downto 4);
                            --FRM_o_B <= C0(to_integer(sv_y_matrix),to_integer(sv_x_matrix))( 3 downto 0);
                        end if;
                        --C1
                        if ((sv_v_cnt >= 120 and sv_v_cnt <= 139 and sv_h_cnt >= 140 and sv_h_cnt <= 199) 
                            or (sv_v_cnt >= 140 and sv_v_cnt <= 159 and sv_h_cnt >= 140 and sv_h_cnt <= 159) 
                            or (sv_v_cnt >= 140 and sv_v_cnt <= 159 and sv_h_cnt >= 180 and sv_h_cnt <= 199) 
                            or (sv_v_cnt >= 160 and sv_v_cnt <= 179 and sv_h_cnt >= 140 and sv_h_cnt <= 199)) then
                            FRM_o_R <= "0000";
                            FRM_o_G <= "0000";
                            FRM_o_B <= "0000";
                        elsif (sv_v_cnt >= 140 and sv_v_cnt <= 159 and sv_h_cnt >= 160 and sv_h_cnt <= 179) then
                            sv_x_matrix <= sv_h_cnt - 160;
                            sv_y_matrix <= sv_v_cnt - 140;
                            if (si_curs_x = 1 and si_curs_y = 2) then
                                st_lamp_off <= C1;
                                FRM_o_R     <= st_cursore(to_integer(sv_y_matrix),to_integer(sv_x_matrix))(11 downto 8);
                                FRM_o_G     <= st_cursore(to_integer(sv_y_matrix),to_integer(sv_x_matrix))( 7 downto 4);
                                FRM_o_B     <= st_cursore(to_integer(sv_y_matrix),to_integer(sv_x_matrix))( 3 downto 0);
                            else
                                FRM_o_R     <= C1(to_integer(sv_y_matrix),to_integer(sv_x_matrix))(11 downto 8);
                                FRM_o_G     <= C1(to_integer(sv_y_matrix),to_integer(sv_x_matrix))( 7 downto 4);
                                FRM_o_B     <= C1(to_integer(sv_y_matrix),to_integer(sv_x_matrix))( 3 downto 0);
                            end if;
                            --FRM_o_R <= C1(to_integer(sv_y_matrix),to_integer(sv_x_matrix))(11 downto 8);
                            --FRM_o_G <= C1(to_integer(sv_y_matrix),to_integer(sv_x_matrix))( 7 downto 4);
                            --FRM_o_B <= C1(to_integer(sv_y_matrix),to_integer(sv_x_matrix))( 3 downto 0);
                        end if;
                        --C2
                        if ((sv_v_cnt >= 120 and sv_v_cnt <= 139 and sv_h_cnt >= 200 and sv_h_cnt <= 259) 
                            or (sv_v_cnt >= 140 and sv_v_cnt <= 159 and sv_h_cnt >= 200 and sv_h_cnt <= 219) 
                            or (sv_v_cnt >= 140 and sv_v_cnt <= 159 and sv_h_cnt >= 240 and sv_h_cnt <= 259) 
                            or (sv_v_cnt >= 160 and sv_v_cnt <= 179 and sv_h_cnt >= 200 and sv_h_cnt <= 259)) then
                            FRM_o_R <= "1111";
                            FRM_o_G <= "1111";
                            FRM_o_B <= "1111";
                        elsif (sv_v_cnt >= 140 and sv_v_cnt <= 159 and sv_h_cnt >= 220 and sv_h_cnt <= 239) then
                            sv_x_matrix <= sv_h_cnt - 220;
                            sv_y_matrix <= sv_v_cnt - 140;
                            if (si_curs_x = 2 and si_curs_y = 2) then
                                st_lamp_off <= C2;
                                FRM_o_R     <= st_cursore(to_integer(sv_y_matrix),to_integer(sv_x_matrix))(11 downto 8);
                                FRM_o_G     <= st_cursore(to_integer(sv_y_matrix),to_integer(sv_x_matrix))( 7 downto 4);
                                FRM_o_B     <= st_cursore(to_integer(sv_y_matrix),to_integer(sv_x_matrix))( 3 downto 0);
                            else
                                FRM_o_R     <= C2(to_integer(sv_y_matrix),to_integer(sv_x_matrix))(11 downto 8);
                                FRM_o_G     <= C2(to_integer(sv_y_matrix),to_integer(sv_x_matrix))( 7 downto 4);
                                FRM_o_B     <= C2(to_integer(sv_y_matrix),to_integer(sv_x_matrix))( 3 downto 0);
                            end if;
                            --FRM_o_R <= C2(to_integer(sv_y_matrix),to_integer(sv_x_matrix))(11 downto 8);
                            --FRM_o_G <= C2(to_integer(sv_y_matrix),to_integer(sv_x_matrix))( 7 downto 4);
                            --FRM_o_B <= C2(to_integer(sv_y_matrix),to_integer(sv_x_matrix))( 3 downto 0);
                        end if;
                        --C3
                        if ((sv_v_cnt >= 120 and sv_v_cnt <= 139 and sv_h_cnt >= 260 and sv_h_cnt <= 319) 
                            or (sv_v_cnt >= 140 and sv_v_cnt <= 159 and sv_h_cnt >= 260 and sv_h_cnt <= 279) 
                            or (sv_v_cnt >= 140 and sv_v_cnt <= 159 and sv_h_cnt >= 300 and sv_h_cnt <= 319) 
                            or (sv_v_cnt >= 160 and sv_v_cnt <= 179 and sv_h_cnt >= 260 and sv_h_cnt <= 319)) then
                            FRM_o_R <= "0000";
                            FRM_o_G <= "0000";
                            FRM_o_B <= "0000";
                        elsif (sv_v_cnt >= 140 and sv_v_cnt <= 159 and sv_h_cnt >= 280 and sv_h_cnt <= 299) then
                            sv_x_matrix <= sv_h_cnt - 280;
                            sv_y_matrix <= sv_v_cnt - 140;
                            if (si_curs_x = 3 and si_curs_y = 2) then
                                st_lamp_off <= C3;
                                FRM_o_R     <= st_cursore(to_integer(sv_y_matrix),to_integer(sv_x_matrix))(11 downto 8);
                                FRM_o_G     <= st_cursore(to_integer(sv_y_matrix),to_integer(sv_x_matrix))( 7 downto 4);
                                FRM_o_B     <= st_cursore(to_integer(sv_y_matrix),to_integer(sv_x_matrix))( 3 downto 0);
                            else
                                FRM_o_R     <= C3(to_integer(sv_y_matrix),to_integer(sv_x_matrix))(11 downto 8);
                                FRM_o_G     <= C3(to_integer(sv_y_matrix),to_integer(sv_x_matrix))( 7 downto 4);
                                FRM_o_B     <= C3(to_integer(sv_y_matrix),to_integer(sv_x_matrix))( 3 downto 0);
                            end if;
                            --FRM_o_R <= C3(to_integer(sv_y_matrix),to_integer(sv_x_matrix))(11 downto 8);
                            --FRM_o_G <= C3(to_integer(sv_y_matrix),to_integer(sv_x_matrix))( 7 downto 4);
                            --FRM_o_B <= C3(to_integer(sv_y_matrix),to_integer(sv_x_matrix))( 3 downto 0);
                        end if;
                        --C4
                        if ((sv_v_cnt >= 120 and sv_v_cnt <= 139 and sv_h_cnt >= 320 and sv_h_cnt <= 379) 
                            or (sv_v_cnt >= 140 and sv_v_cnt <= 159 and sv_h_cnt >= 320 and sv_h_cnt <= 339) 
                            or (sv_v_cnt >= 140 and sv_v_cnt <= 159 and sv_h_cnt >= 360 and sv_h_cnt <= 379) 
                            or (sv_v_cnt >= 160 and sv_v_cnt <= 179 and sv_h_cnt >= 320 and sv_h_cnt <= 379)) then
                            FRM_o_R <= "1111";
                            FRM_o_G <= "1111";
                            FRM_o_B <= "1111";
                        elsif (sv_v_cnt >= 140 and sv_v_cnt <= 159 and sv_h_cnt >= 340 and sv_h_cnt <= 359) then
                            sv_x_matrix <= sv_h_cnt - 340;
                            sv_y_matrix <= sv_v_cnt - 140;
                            if (si_curs_x = 4 and si_curs_y = 2) then
                                st_lamp_off <= C4;
                                FRM_o_R     <= st_cursore(to_integer(sv_y_matrix),to_integer(sv_x_matrix))(11 downto 8);
                                FRM_o_G     <= st_cursore(to_integer(sv_y_matrix),to_integer(sv_x_matrix))( 7 downto 4);
                                FRM_o_B     <= st_cursore(to_integer(sv_y_matrix),to_integer(sv_x_matrix))( 3 downto 0);
                            else
                                FRM_o_R     <= C4(to_integer(sv_y_matrix),to_integer(sv_x_matrix))(11 downto 8);
                                FRM_o_G     <= C4(to_integer(sv_y_matrix),to_integer(sv_x_matrix))( 7 downto 4);
                                FRM_o_B     <= C4(to_integer(sv_y_matrix),to_integer(sv_x_matrix))( 3 downto 0);
                            end if;
                            --FRM_o_R <= C4(to_integer(sv_y_matrix),to_integer(sv_x_matrix))(11 downto 8);
                            --FRM_o_G <= C4(to_integer(sv_y_matrix),to_integer(sv_x_matrix))( 7 downto 4);
                            --FRM_o_B <= C4(to_integer(sv_y_matrix),to_integer(sv_x_matrix))( 3 downto 0);
                        end if;
                        --C5
                        if ((sv_v_cnt >= 120 and sv_v_cnt <= 139 and sv_h_cnt >= 380 and sv_h_cnt <= 439) 
                            or (sv_v_cnt >= 140 and sv_v_cnt <= 159 and sv_h_cnt >= 380 and sv_h_cnt <= 399) 
                            or (sv_v_cnt >= 140 and sv_v_cnt <= 159 and sv_h_cnt >= 420 and sv_h_cnt <= 439) 
                            or (sv_v_cnt >= 160 and sv_v_cnt <= 179 and sv_h_cnt >= 380 and sv_h_cnt <= 439)) then
                            FRM_o_R <= "0000";
                            FRM_o_G <= "0000";
                            FRM_o_B <= "0000";
                        elsif (sv_v_cnt >= 140 and sv_v_cnt <= 159 and sv_h_cnt >= 400 and sv_h_cnt <= 419) then
                            sv_x_matrix <= sv_h_cnt - 400;
                            sv_y_matrix <= sv_v_cnt - 140;
                            if (si_curs_x = 5 and si_curs_y = 2) then
                                st_lamp_off <= C5;
                                FRM_o_R     <= st_cursore(to_integer(sv_y_matrix),to_integer(sv_x_matrix))(11 downto 8);
                                FRM_o_G     <= st_cursore(to_integer(sv_y_matrix),to_integer(sv_x_matrix))( 7 downto 4);
                                FRM_o_B     <= st_cursore(to_integer(sv_y_matrix),to_integer(sv_x_matrix))( 3 downto 0);
                            else
                                FRM_o_R     <= C5(to_integer(sv_y_matrix),to_integer(sv_x_matrix))(11 downto 8);
                                FRM_o_G     <= C5(to_integer(sv_y_matrix),to_integer(sv_x_matrix))( 7 downto 4);
                                FRM_o_B     <= C5(to_integer(sv_y_matrix),to_integer(sv_x_matrix))( 3 downto 0);
                            end if;
                            --FRM_o_R <= C5(to_integer(sv_y_matrix),to_integer(sv_x_matrix))(11 downto 8);
                            --FRM_o_G <= C5(to_integer(sv_y_matrix),to_integer(sv_x_matrix))( 7 downto 4);
                            --FRM_o_B <= C5(to_integer(sv_y_matrix),to_integer(sv_x_matrix))( 3 downto 0);
                        end if;
                        --C6
                        if ((sv_v_cnt >= 120 and sv_v_cnt <= 139 and sv_h_cnt >= 440 and sv_h_cnt <= 499) 
                            or (sv_v_cnt >= 140 and sv_v_cnt <= 159 and sv_h_cnt >= 440 and sv_h_cnt <= 459) 
                            or (sv_v_cnt >= 140 and sv_v_cnt <= 159 and sv_h_cnt >= 480 and sv_h_cnt <= 499) 
                            or (sv_v_cnt >= 160 and sv_v_cnt <= 179 and sv_h_cnt >= 440 and sv_h_cnt <= 499)) then
                            FRM_o_R <= "1111";
                            FRM_o_G <= "1111";
                            FRM_o_B <= "1111";
                        elsif (sv_v_cnt >= 140 and sv_v_cnt <= 159 and sv_h_cnt >= 460 and sv_h_cnt <= 479) then
                            sv_x_matrix <= sv_h_cnt - 460;
                            sv_y_matrix <= sv_v_cnt - 140;
                            if (si_curs_x = 6 and si_curs_y = 2) then
                                st_lamp_off <= C6;
                                FRM_o_R     <= st_cursore(to_integer(sv_y_matrix),to_integer(sv_x_matrix))(11 downto 8);
                                FRM_o_G     <= st_cursore(to_integer(sv_y_matrix),to_integer(sv_x_matrix))( 7 downto 4);
                                FRM_o_B     <= st_cursore(to_integer(sv_y_matrix),to_integer(sv_x_matrix))( 3 downto 0);
                            else
                                FRM_o_R     <= C6(to_integer(sv_y_matrix),to_integer(sv_x_matrix))(11 downto 8);
                                FRM_o_G     <= C6(to_integer(sv_y_matrix),to_integer(sv_x_matrix))( 7 downto 4);
                                FRM_o_B     <= C6(to_integer(sv_y_matrix),to_integer(sv_x_matrix))( 3 downto 0);
                            end if;
                            --FRM_o_R <= C6(to_integer(sv_y_matrix),to_integer(sv_x_matrix))(11 downto 8);
                            --FRM_o_G <= C6(to_integer(sv_y_matrix),to_integer(sv_x_matrix))( 7 downto 4);
                            --FRM_o_B <= C6(to_integer(sv_y_matrix),to_integer(sv_x_matrix))( 3 downto 0);
                        end if;
                        --C7
                        if ((sv_v_cnt >= 120 and sv_v_cnt <= 139 and sv_h_cnt >= 500 and sv_h_cnt <= 559) 
                            or (sv_v_cnt >= 140 and sv_v_cnt <= 159 and sv_h_cnt >= 500 and sv_h_cnt <= 519) 
                            or (sv_v_cnt >= 140 and sv_v_cnt <= 159 and sv_h_cnt >= 540 and sv_h_cnt <= 559) 
                            or (sv_v_cnt >= 160 and sv_v_cnt <= 179 and sv_h_cnt >= 500 and sv_h_cnt <= 559)) then
                            FRM_o_R <= "0000";
                            FRM_o_G <= "0000";
                            FRM_o_B <= "0000";
                        elsif (sv_v_cnt >= 140 and sv_v_cnt <= 159 and sv_h_cnt >= 520 and sv_h_cnt <= 539) then
                            sv_x_matrix <= sv_h_cnt - 520;
                            sv_y_matrix <= sv_v_cnt - 140;
                            if (si_curs_x = 7 and si_curs_y = 2) then
                                st_lamp_off <= C7;
                                FRM_o_R     <= st_cursore(to_integer(sv_y_matrix),to_integer(sv_x_matrix))(11 downto 8);
                                FRM_o_G     <= st_cursore(to_integer(sv_y_matrix),to_integer(sv_x_matrix))( 7 downto 4);
                                FRM_o_B     <= st_cursore(to_integer(sv_y_matrix),to_integer(sv_x_matrix))( 3 downto 0);
                            else
                                FRM_o_R     <= C7(to_integer(sv_y_matrix),to_integer(sv_x_matrix))(11 downto 8);
                                FRM_o_G     <= C7(to_integer(sv_y_matrix),to_integer(sv_x_matrix))( 7 downto 4);
                                FRM_o_B     <= C7(to_integer(sv_y_matrix),to_integer(sv_x_matrix))( 3 downto 0);
                            end if;
                            --FRM_o_R <= C7(to_integer(sv_y_matrix),to_integer(sv_x_matrix))(11 downto 8);
                            --FRM_o_G <= C7(to_integer(sv_y_matrix),to_integer(sv_x_matrix))( 7 downto 4);
                            --FRM_o_B <= C7(to_integer(sv_y_matrix),to_integer(sv_x_matrix))( 3 downto 0);
                        end if;
                        --D0
                        if ((sv_v_cnt >= 180 and sv_v_cnt <= 199 and sv_h_cnt >= 80 and sv_h_cnt <= 139) 
                            or (sv_v_cnt >= 200 and sv_v_cnt <= 219 and sv_h_cnt >= 80 and sv_h_cnt <= 99) 
                            or (sv_v_cnt >= 200 and sv_v_cnt <= 219 and sv_h_cnt >= 120 and sv_h_cnt <= 139) 
                            or (sv_v_cnt >= 220 and sv_v_cnt <= 239 and sv_h_cnt >= 80 and sv_h_cnt <= 139)) then
                            FRM_o_R <= "0000";
                            FRM_o_G <= "0000";
                            FRM_o_B <= "0000";
                        elsif (sv_v_cnt >= 200 and sv_v_cnt <= 219 and sv_h_cnt >= 100 and sv_h_cnt <= 119) then
                            sv_x_matrix <= sv_h_cnt - 100;
                            sv_y_matrix <= sv_v_cnt - 200;
                            if (si_curs_x = 0 and si_curs_y = 3) then
                                st_lamp_off <= D0;
                                FRM_o_R     <= st_cursore(to_integer(sv_y_matrix),to_integer(sv_x_matrix))(11 downto 8);
                                FRM_o_G     <= st_cursore(to_integer(sv_y_matrix),to_integer(sv_x_matrix))( 7 downto 4);
                                FRM_o_B     <= st_cursore(to_integer(sv_y_matrix),to_integer(sv_x_matrix))( 3 downto 0);
                            else
                                FRM_o_R     <= D0(to_integer(sv_y_matrix),to_integer(sv_x_matrix))(11 downto 8);
                                FRM_o_G     <= D0(to_integer(sv_y_matrix),to_integer(sv_x_matrix))( 7 downto 4);
                                FRM_o_B     <= D0(to_integer(sv_y_matrix),to_integer(sv_x_matrix))( 3 downto 0);
                            end if;
                            --FRM_o_R <= D0(to_integer(sv_y_matrix),to_integer(sv_x_matrix))(11 downto 8);
                            --FRM_o_G <= D0(to_integer(sv_y_matrix),to_integer(sv_x_matrix))( 7 downto 4);
                            --FRM_o_B <= D0(to_integer(sv_y_matrix),to_integer(sv_x_matrix))( 3 downto 0);
                        end if;
                        --D1
                        if ((sv_v_cnt >= 180 and sv_v_cnt <= 199 and sv_h_cnt >= 140 and sv_h_cnt <= 199) 
                            or (sv_v_cnt >= 200 and sv_v_cnt <= 219 and sv_h_cnt >= 140 and sv_h_cnt <= 159) 
                            or (sv_v_cnt >= 200 and sv_v_cnt <= 219 and sv_h_cnt >= 180 and sv_h_cnt <= 199) 
                            or (sv_v_cnt >= 220 and sv_v_cnt <= 239 and sv_h_cnt >= 140 and sv_h_cnt <= 199)) then
                            FRM_o_R <= "1111";
                            FRM_o_G <= "1111";
                            FRM_o_B <= "1111";
                        elsif (sv_v_cnt >= 200 and sv_v_cnt <= 219 and sv_h_cnt >= 160 and sv_h_cnt <= 179) then
                            sv_x_matrix <= sv_h_cnt - 160;
                            sv_y_matrix <= sv_v_cnt - 200;
                            if (si_curs_x = 1 and si_curs_y = 3) then
                                st_lamp_off <= D1;
                                FRM_o_R     <= st_cursore(to_integer(sv_y_matrix),to_integer(sv_x_matrix))(11 downto 8);
                                FRM_o_G     <= st_cursore(to_integer(sv_y_matrix),to_integer(sv_x_matrix))( 7 downto 4);
                                FRM_o_B     <= st_cursore(to_integer(sv_y_matrix),to_integer(sv_x_matrix))( 3 downto 0);
                            else
                                FRM_o_R     <= D1(to_integer(sv_y_matrix),to_integer(sv_x_matrix))(11 downto 8);
                                FRM_o_G     <= D1(to_integer(sv_y_matrix),to_integer(sv_x_matrix))( 7 downto 4);
                                FRM_o_B     <= D1(to_integer(sv_y_matrix),to_integer(sv_x_matrix))( 3 downto 0);
                            end if;
                            --FRM_o_R <= D1(to_integer(sv_y_matrix),to_integer(sv_x_matrix))(11 downto 8);
                            --FRM_o_G <= D1(to_integer(sv_y_matrix),to_integer(sv_x_matrix))( 7 downto 4);
                            --FRM_o_B <= D1(to_integer(sv_y_matrix),to_integer(sv_x_matrix))( 3 downto 0);
                        end if;
                        --D2
                        if ((sv_v_cnt >= 180 and sv_v_cnt <= 199 and sv_h_cnt >= 200 and sv_h_cnt <= 259) 
                            or (sv_v_cnt >= 200 and sv_v_cnt <= 219 and sv_h_cnt >= 200 and sv_h_cnt <= 219) 
                            or (sv_v_cnt >= 200 and sv_v_cnt <= 219 and sv_h_cnt >= 240 and sv_h_cnt <= 259) 
                            or (sv_v_cnt >= 220 and sv_v_cnt <= 239 and sv_h_cnt >= 200 and sv_h_cnt <= 259)) then
                            FRM_o_R <= "0000";
                            FRM_o_G <= "0000";
                            FRM_o_B <= "0000";
                        elsif (sv_v_cnt >= 200 and sv_v_cnt <= 219 and sv_h_cnt >= 220 and sv_h_cnt <= 239) then
                            sv_x_matrix <= sv_h_cnt - 220;
                            sv_y_matrix <= sv_v_cnt - 200;
                            if (si_curs_x = 2 and si_curs_y = 3) then
                                st_lamp_off <= D2;
                                FRM_o_R     <= st_cursore(to_integer(sv_y_matrix),to_integer(sv_x_matrix))(11 downto 8);
                                FRM_o_G     <= st_cursore(to_integer(sv_y_matrix),to_integer(sv_x_matrix))( 7 downto 4);
                                FRM_o_B     <= st_cursore(to_integer(sv_y_matrix),to_integer(sv_x_matrix))( 3 downto 0);
                            else
                                FRM_o_R     <= D2(to_integer(sv_y_matrix),to_integer(sv_x_matrix))(11 downto 8);
                                FRM_o_G     <= D2(to_integer(sv_y_matrix),to_integer(sv_x_matrix))( 7 downto 4);
                                FRM_o_B     <= D2(to_integer(sv_y_matrix),to_integer(sv_x_matrix))( 3 downto 0);
                            end if;
                            --FRM_o_R <= D2(to_integer(sv_y_matrix),to_integer(sv_x_matrix))(11 downto 8);
                            --FRM_o_G <= D2(to_integer(sv_y_matrix),to_integer(sv_x_matrix))( 7 downto 4);
                            --FRM_o_B <= D2(to_integer(sv_y_matrix),to_integer(sv_x_matrix))( 3 downto 0);
                        end if;
                        --D3
                        if ((sv_v_cnt >= 180 and sv_v_cnt <= 199 and sv_h_cnt >= 260 and sv_h_cnt <= 319) 
                            or (sv_v_cnt >= 200 and sv_v_cnt <= 219 and sv_h_cnt >= 260 and sv_h_cnt <= 279) 
                            or (sv_v_cnt >= 200 and sv_v_cnt <= 219 and sv_h_cnt >= 300 and sv_h_cnt <= 319) 
                            or (sv_v_cnt >= 220 and sv_v_cnt <= 239 and sv_h_cnt >= 260 and sv_h_cnt <= 319)) then
                            FRM_o_R <= "1111";
                            FRM_o_G <= "1111";
                            FRM_o_B <= "1111";
                        elsif (sv_v_cnt >= 200 and sv_v_cnt <= 219 and sv_h_cnt >= 280 and sv_h_cnt <= 299) then
                            sv_x_matrix <= sv_h_cnt - 280;
                            sv_y_matrix <= sv_v_cnt - 200;
                            if (si_curs_x = 3 and si_curs_y = 3) then
                                st_lamp_off <= D3;
                                FRM_o_R     <= st_cursore(to_integer(sv_y_matrix),to_integer(sv_x_matrix))(11 downto 8);
                                FRM_o_G     <= st_cursore(to_integer(sv_y_matrix),to_integer(sv_x_matrix))( 7 downto 4);
                                FRM_o_B     <= st_cursore(to_integer(sv_y_matrix),to_integer(sv_x_matrix))( 3 downto 0);
                            else
                                FRM_o_R     <= D3(to_integer(sv_y_matrix),to_integer(sv_x_matrix))(11 downto 8);
                                FRM_o_G     <= D3(to_integer(sv_y_matrix),to_integer(sv_x_matrix))( 7 downto 4);
                                FRM_o_B     <= D3(to_integer(sv_y_matrix),to_integer(sv_x_matrix))( 3 downto 0);
                            end if;
                            --FRM_o_R <= D3(to_integer(sv_y_matrix),to_integer(sv_x_matrix))(11 downto 8);
                            --FRM_o_G <= D3(to_integer(sv_y_matrix),to_integer(sv_x_matrix))( 7 downto 4);
                            --FRM_o_B <= D3(to_integer(sv_y_matrix),to_integer(sv_x_matrix))( 3 downto 0);
                        end if;
                        --D4
                        if ((sv_v_cnt >= 180 and sv_v_cnt <= 199 and sv_h_cnt >= 320 and sv_h_cnt <= 379) 
                            or (sv_v_cnt >= 200 and sv_v_cnt <= 219 and sv_h_cnt >= 320 and sv_h_cnt <= 339) 
                            or (sv_v_cnt >= 200 and sv_v_cnt <= 219 and sv_h_cnt >= 360 and sv_h_cnt <= 379) 
                            or (sv_v_cnt >= 220 and sv_v_cnt <= 239 and sv_h_cnt >= 320 and sv_h_cnt <= 379)) then
                            FRM_o_R <= "0000";
                            FRM_o_G <= "0000";
                            FRM_o_B <= "0000";
                        elsif (sv_v_cnt >= 200 and sv_v_cnt <= 219 and sv_h_cnt >= 340 and sv_h_cnt <= 359) then
                            sv_x_matrix <= sv_h_cnt - 340;
                            sv_y_matrix <= sv_v_cnt - 200;
                            if (si_curs_x = 4 and si_curs_y = 3) then
                                st_lamp_off <= D4;
                                FRM_o_R     <= st_cursore(to_integer(sv_y_matrix),to_integer(sv_x_matrix))(11 downto 8);
                                FRM_o_G     <= st_cursore(to_integer(sv_y_matrix),to_integer(sv_x_matrix))( 7 downto 4);
                                FRM_o_B     <= st_cursore(to_integer(sv_y_matrix),to_integer(sv_x_matrix))( 3 downto 0);
                            else
                                FRM_o_R     <= D4(to_integer(sv_y_matrix),to_integer(sv_x_matrix))(11 downto 8);
                                FRM_o_G     <= D4(to_integer(sv_y_matrix),to_integer(sv_x_matrix))( 7 downto 4);
                                FRM_o_B     <= D4(to_integer(sv_y_matrix),to_integer(sv_x_matrix))( 3 downto 0);
                            end if;
                            --FRM_o_R <= D4(to_integer(sv_y_matrix),to_integer(sv_x_matrix))(11 downto 8);
                            --FRM_o_G <= D4(to_integer(sv_y_matrix),to_integer(sv_x_matrix))( 7 downto 4);
                            --FRM_o_B <= D4(to_integer(sv_y_matrix),to_integer(sv_x_matrix))( 3 downto 0);
                        end if;
                        --D5
                        if ((sv_v_cnt >= 180 and sv_v_cnt <= 199 and sv_h_cnt >= 380 and sv_h_cnt <= 439) 
                            or (sv_v_cnt >= 200 and sv_v_cnt <= 219 and sv_h_cnt >= 380 and sv_h_cnt <= 399) 
                            or (sv_v_cnt >= 200 and sv_v_cnt <= 219 and sv_h_cnt >= 420 and sv_h_cnt <= 439) 
                            or (sv_v_cnt >= 220 and sv_v_cnt <= 239 and sv_h_cnt >= 380 and sv_h_cnt <= 439)) then
                            FRM_o_R <= "1111";
                            FRM_o_G <= "1111";
                            FRM_o_B <= "1111";
                        elsif (sv_v_cnt >= 200 and sv_v_cnt <= 219 and sv_h_cnt >= 400 and sv_h_cnt <= 419) then
                            sv_x_matrix <= sv_h_cnt - 400;
                            sv_y_matrix <= sv_v_cnt - 200;
                            if (si_curs_x = 5 and si_curs_y = 3) then
                                st_lamp_off <= D5;
                                FRM_o_R     <= st_cursore(to_integer(sv_y_matrix),to_integer(sv_x_matrix))(11 downto 8);
                                FRM_o_G     <= st_cursore(to_integer(sv_y_matrix),to_integer(sv_x_matrix))( 7 downto 4);
                                FRM_o_B     <= st_cursore(to_integer(sv_y_matrix),to_integer(sv_x_matrix))( 3 downto 0);
                            else
                                FRM_o_R     <= D5(to_integer(sv_y_matrix),to_integer(sv_x_matrix))(11 downto 8);
                                FRM_o_G     <= D5(to_integer(sv_y_matrix),to_integer(sv_x_matrix))( 7 downto 4);
                                FRM_o_B     <= D5(to_integer(sv_y_matrix),to_integer(sv_x_matrix))( 3 downto 0);
                            end if;
                            --FRM_o_R <= D5(to_integer(sv_y_matrix),to_integer(sv_x_matrix))(11 downto 8);
                            --FRM_o_G <= D5(to_integer(sv_y_matrix),to_integer(sv_x_matrix))( 7 downto 4);
                            --FRM_o_B <= D5(to_integer(sv_y_matrix),to_integer(sv_x_matrix))( 3 downto 0);
                        end if;
                        --D6
                        if ((sv_v_cnt >= 180 and sv_v_cnt <= 199 and sv_h_cnt >= 440 and sv_h_cnt <= 499) 
                            or (sv_v_cnt >= 200 and sv_v_cnt <= 219 and sv_h_cnt >= 440 and sv_h_cnt <= 459) 
                            or (sv_v_cnt >= 200 and sv_v_cnt <= 219 and sv_h_cnt >= 480 and sv_h_cnt <= 499) 
                            or (sv_v_cnt >= 220 and sv_v_cnt <= 239 and sv_h_cnt >= 440 and sv_h_cnt <= 499)) then
                            FRM_o_R <= "0000";
                            FRM_o_G <= "0000";
                            FRM_o_B <= "0000";
                        elsif (sv_v_cnt >= 200 and sv_v_cnt <= 219 and sv_h_cnt >= 460 and sv_h_cnt <= 479) then
                            sv_x_matrix <= sv_h_cnt - 460;
                            sv_y_matrix <= sv_v_cnt - 200;
                            if (si_curs_x = 6 and si_curs_y = 3) then
                                st_lamp_off <= D6;
                                FRM_o_R     <= st_cursore(to_integer(sv_y_matrix),to_integer(sv_x_matrix))(11 downto 8);
                                FRM_o_G     <= st_cursore(to_integer(sv_y_matrix),to_integer(sv_x_matrix))( 7 downto 4);
                                FRM_o_B     <= st_cursore(to_integer(sv_y_matrix),to_integer(sv_x_matrix))( 3 downto 0);
                            else
                                FRM_o_R     <= D6(to_integer(sv_y_matrix),to_integer(sv_x_matrix))(11 downto 8);
                                FRM_o_G     <= D6(to_integer(sv_y_matrix),to_integer(sv_x_matrix))( 7 downto 4);
                                FRM_o_B     <= D6(to_integer(sv_y_matrix),to_integer(sv_x_matrix))( 3 downto 0);
                            end if;
                            --FRM_o_R <= D6(to_integer(sv_y_matrix),to_integer(sv_x_matrix))(11 downto 8);
                            --FRM_o_G <= D6(to_integer(sv_y_matrix),to_integer(sv_x_matrix))( 7 downto 4);
                            --FRM_o_B <= D6(to_integer(sv_y_matrix),to_integer(sv_x_matrix))( 3 downto 0);
                        end if;
                        --D7
                        if ((sv_v_cnt >= 180 and sv_v_cnt <= 199 and sv_h_cnt >= 500 and sv_h_cnt <= 559) 
                            or (sv_v_cnt >= 200 and sv_v_cnt <= 219 and sv_h_cnt >= 500 and sv_h_cnt <= 519) 
                            or (sv_v_cnt >= 200 and sv_v_cnt <= 219 and sv_h_cnt >= 540 and sv_h_cnt <= 559) 
                            or (sv_v_cnt >= 220 and sv_v_cnt <= 239 and sv_h_cnt >= 500 and sv_h_cnt <= 559)) then
                            FRM_o_R <= "1111";
                            FRM_o_G <= "1111";
                            FRM_o_B <= "1111";
                        elsif (sv_v_cnt >= 200 and sv_v_cnt <= 219 and sv_h_cnt >= 520 and sv_h_cnt <= 539) then
                            sv_x_matrix <= sv_h_cnt - 520;
                            sv_y_matrix <= sv_v_cnt - 200;
                            if (si_curs_x = 7 and si_curs_y = 3) then
                                st_lamp_off <= D7;
                                FRM_o_R     <= st_cursore(to_integer(sv_y_matrix),to_integer(sv_x_matrix))(11 downto 8);
                                FRM_o_G     <= st_cursore(to_integer(sv_y_matrix),to_integer(sv_x_matrix))( 7 downto 4);
                                FRM_o_B     <= st_cursore(to_integer(sv_y_matrix),to_integer(sv_x_matrix))( 3 downto 0);
                            else
                                FRM_o_R     <= D7(to_integer(sv_y_matrix),to_integer(sv_x_matrix))(11 downto 8);
                                FRM_o_G     <= D7(to_integer(sv_y_matrix),to_integer(sv_x_matrix))( 7 downto 4);
                                FRM_o_B     <= D7(to_integer(sv_y_matrix),to_integer(sv_x_matrix))( 3 downto 0);
                            end if;
                            --FRM_o_R <= D7(to_integer(sv_y_matrix),to_integer(sv_x_matrix))(11 downto 8);
                            --FRM_o_G <= D7(to_integer(sv_y_matrix),to_integer(sv_x_matrix))( 7 downto 4);
                            --FRM_o_B <= D7(to_integer(sv_y_matrix),to_integer(sv_x_matrix))( 3 downto 0);
                        end if;
                        --E0
                        if ((sv_v_cnt >= 240 and sv_v_cnt <= 259 and sv_h_cnt >= 80 and sv_h_cnt <= 139) 
                            or (sv_v_cnt >= 260 and sv_v_cnt <= 279 and sv_h_cnt >= 80 and sv_h_cnt <= 99) 
                            or (sv_v_cnt >= 260 and sv_v_cnt <= 279 and sv_h_cnt >= 120 and sv_h_cnt <= 139) 
                            or (sv_v_cnt >= 280 and sv_v_cnt <= 299 and sv_h_cnt >= 80 and sv_h_cnt <= 139)) then
                            FRM_o_R <= "1111";
                            FRM_o_G <= "1111";
                            FRM_o_B <= "1111";
                        elsif (sv_v_cnt >= 260 and sv_v_cnt <= 279 and sv_h_cnt >= 100 and sv_h_cnt <= 119) then
                            sv_x_matrix <= sv_h_cnt - 100;
                            sv_y_matrix <= sv_v_cnt - 260;
                            if (si_curs_x = 0 and si_curs_y = 4) then
                                st_lamp_off <= E0;
                                FRM_o_R     <= st_cursore(to_integer(sv_y_matrix),to_integer(sv_x_matrix))(11 downto 8);
                                FRM_o_G     <= st_cursore(to_integer(sv_y_matrix),to_integer(sv_x_matrix))( 7 downto 4);
                                FRM_o_B     <= st_cursore(to_integer(sv_y_matrix),to_integer(sv_x_matrix))( 3 downto 0);
                            else
                                FRM_o_R     <= E0(to_integer(sv_y_matrix),to_integer(sv_x_matrix))(11 downto 8);
                                FRM_o_G     <= E0(to_integer(sv_y_matrix),to_integer(sv_x_matrix))( 7 downto 4);
                                FRM_o_B     <= E0(to_integer(sv_y_matrix),to_integer(sv_x_matrix))( 3 downto 0);
                            end if;
                            --FRM_o_R <= E0(to_integer(sv_y_matrix),to_integer(sv_x_matrix))(11 downto 8);
                            --FRM_o_G <= E0(to_integer(sv_y_matrix),to_integer(sv_x_matrix))( 7 downto 4);
                            --FRM_o_B <= E0(to_integer(sv_y_matrix),to_integer(sv_x_matrix))( 3 downto 0);
                        end if;
                        --E1
                        if ((sv_v_cnt >= 240 and sv_v_cnt <= 259 and sv_h_cnt >= 140 and sv_h_cnt <= 199) 
                            or (sv_v_cnt >= 260 and sv_v_cnt <= 279 and sv_h_cnt >= 140 and sv_h_cnt <= 159) 
                            or (sv_v_cnt >= 260 and sv_v_cnt <= 279 and sv_h_cnt >= 180 and sv_h_cnt <= 199) 
                            or (sv_v_cnt >= 280 and sv_v_cnt <= 299 and sv_h_cnt >= 140 and sv_h_cnt <= 199)) then
                            FRM_o_R <= "0000";
                            FRM_o_G <= "0000";
                            FRM_o_B <= "0000";
                        elsif (sv_v_cnt >= 260 and sv_v_cnt <= 279 and sv_h_cnt >= 160 and sv_h_cnt <= 179) then
                            sv_x_matrix <= sv_h_cnt - 160;
                            sv_y_matrix <= sv_v_cnt - 260;
                            if (si_curs_x = 1 and si_curs_y = 4) then
                                st_lamp_off <= E1;
                                FRM_o_R     <= st_cursore(to_integer(sv_y_matrix),to_integer(sv_x_matrix))(11 downto 8);
                                FRM_o_G     <= st_cursore(to_integer(sv_y_matrix),to_integer(sv_x_matrix))( 7 downto 4);
                                FRM_o_B     <= st_cursore(to_integer(sv_y_matrix),to_integer(sv_x_matrix))( 3 downto 0);
                            else
                                FRM_o_R     <= E1(to_integer(sv_y_matrix),to_integer(sv_x_matrix))(11 downto 8);
                                FRM_o_G     <= E1(to_integer(sv_y_matrix),to_integer(sv_x_matrix))( 7 downto 4);
                                FRM_o_B     <= E1(to_integer(sv_y_matrix),to_integer(sv_x_matrix))( 3 downto 0);
                            end if;
                            --FRM_o_R <= E1(to_integer(sv_y_matrix),to_integer(sv_x_matrix))(11 downto 8);
                            --FRM_o_G <= E1(to_integer(sv_y_matrix),to_integer(sv_x_matrix))( 7 downto 4);
                            --FRM_o_B <= E1(to_integer(sv_y_matrix),to_integer(sv_x_matrix))( 3 downto 0);
                        end if;
                        --E2
                        if ((sv_v_cnt >= 240 and sv_v_cnt <= 259 and sv_h_cnt >= 200 and sv_h_cnt <= 259) 
                            or (sv_v_cnt >= 260 and sv_v_cnt <= 279 and sv_h_cnt >= 200 and sv_h_cnt <= 219) 
                            or (sv_v_cnt >= 260 and sv_v_cnt <= 279 and sv_h_cnt >= 240 and sv_h_cnt <= 259) 
                            or (sv_v_cnt >= 280 and sv_v_cnt <= 299 and sv_h_cnt >= 200 and sv_h_cnt <= 259)) then
                            FRM_o_R <= "1111";
                            FRM_o_G <= "1111";
                            FRM_o_B <= "1111";
                        elsif (sv_v_cnt >= 260 and sv_v_cnt <= 279 and sv_h_cnt >= 220 and sv_h_cnt <= 239) then
                            sv_x_matrix <= sv_h_cnt - 220;
                            sv_y_matrix <= sv_v_cnt - 260;
                            if (si_curs_x = 2 and si_curs_y = 4) then
                                st_lamp_off <= E2;
                                FRM_o_R     <= st_cursore(to_integer(sv_y_matrix),to_integer(sv_x_matrix))(11 downto 8);
                                FRM_o_G     <= st_cursore(to_integer(sv_y_matrix),to_integer(sv_x_matrix))( 7 downto 4);
                                FRM_o_B     <= st_cursore(to_integer(sv_y_matrix),to_integer(sv_x_matrix))( 3 downto 0);
                            else
                                FRM_o_R     <= E2(to_integer(sv_y_matrix),to_integer(sv_x_matrix))(11 downto 8);
                                FRM_o_G     <= E2(to_integer(sv_y_matrix),to_integer(sv_x_matrix))( 7 downto 4);
                                FRM_o_B     <= E2(to_integer(sv_y_matrix),to_integer(sv_x_matrix))( 3 downto 0);
                            end if;
                            --RM_o_R <= E2(to_integer(sv_y_matrix),to_integer(sv_x_matrix))(11 downto 8);
                            --RM_o_G <= E2(to_integer(sv_y_matrix),to_integer(sv_x_matrix))( 7 downto 4);
                            --RM_o_B <= E2(to_integer(sv_y_matrix),to_integer(sv_x_matrix))( 3 downto 0);
                        end if;
                        --E3
                        if ((sv_v_cnt >= 240 and sv_v_cnt <= 259 and sv_h_cnt >= 260 and sv_h_cnt <= 319) 
                            or (sv_v_cnt >= 260 and sv_v_cnt <= 279 and sv_h_cnt >= 260 and sv_h_cnt <= 279) 
                            or (sv_v_cnt >= 260 and sv_v_cnt <= 279 and sv_h_cnt >= 300 and sv_h_cnt <= 319) 
                            or (sv_v_cnt >= 280 and sv_v_cnt <= 299 and sv_h_cnt >= 260 and sv_h_cnt <= 319)) then
                            FRM_o_R <= "0000";
                            FRM_o_G <= "0000";
                            FRM_o_B <= "0000";
                        elsif (sv_v_cnt >= 260 and sv_v_cnt <= 279 and sv_h_cnt >= 280 and sv_h_cnt <= 299) then
                            sv_x_matrix <= sv_h_cnt - 280;
                            sv_y_matrix <= sv_v_cnt - 260;
                            if (si_curs_x = 3 and si_curs_y = 4) then
                                st_lamp_off <= E3;
                                FRM_o_R     <= st_cursore(to_integer(sv_y_matrix),to_integer(sv_x_matrix))(11 downto 8);
                                FRM_o_G     <= st_cursore(to_integer(sv_y_matrix),to_integer(sv_x_matrix))( 7 downto 4);
                                FRM_o_B     <= st_cursore(to_integer(sv_y_matrix),to_integer(sv_x_matrix))( 3 downto 0);
                            else
                                FRM_o_R     <= E3(to_integer(sv_y_matrix),to_integer(sv_x_matrix))(11 downto 8);
                                FRM_o_G     <= E3(to_integer(sv_y_matrix),to_integer(sv_x_matrix))( 7 downto 4);
                                FRM_o_B     <= E3(to_integer(sv_y_matrix),to_integer(sv_x_matrix))( 3 downto 0);
                            end if;
                            --FRM_o_R <= E3(to_integer(sv_y_matrix),to_integer(sv_x_matrix))(11 downto 8);
                            --FRM_o_G <= E3(to_integer(sv_y_matrix),to_integer(sv_x_matrix))( 7 downto 4);
                            --FRM_o_B <= E3(to_integer(sv_y_matrix),to_integer(sv_x_matrix))( 3 downto 0);
                        end if;
                        --E4
                        if ((sv_v_cnt >= 240 and sv_v_cnt <= 259 and sv_h_cnt >= 320 and sv_h_cnt <= 379) 
                            or (sv_v_cnt >= 260 and sv_v_cnt <= 279 and sv_h_cnt >= 320 and sv_h_cnt <= 339) 
                            or (sv_v_cnt >= 260 and sv_v_cnt <= 279 and sv_h_cnt >= 360 and sv_h_cnt <= 379) 
                            or (sv_v_cnt >= 280 and sv_v_cnt <= 299 and sv_h_cnt >= 320 and sv_h_cnt <= 379)) then
                            FRM_o_R <= "1111";
                            FRM_o_G <= "1111";
                            FRM_o_B <= "1111";
                        elsif (sv_v_cnt >= 260 and sv_v_cnt <= 279 and sv_h_cnt >= 340 and sv_h_cnt <= 359) then
                            sv_x_matrix <= sv_h_cnt - 340;
                            sv_y_matrix <= sv_v_cnt - 260;
                            if (si_curs_x = 4 and si_curs_y = 4) then
                                st_lamp_off <= E4;
                                FRM_o_R     <= st_cursore(to_integer(sv_y_matrix),to_integer(sv_x_matrix))(11 downto 8);
                                FRM_o_G     <= st_cursore(to_integer(sv_y_matrix),to_integer(sv_x_matrix))( 7 downto 4);
                                FRM_o_B     <= st_cursore(to_integer(sv_y_matrix),to_integer(sv_x_matrix))( 3 downto 0);
                            else
                                FRM_o_R     <= E4(to_integer(sv_y_matrix),to_integer(sv_x_matrix))(11 downto 8);
                                FRM_o_G     <= E4(to_integer(sv_y_matrix),to_integer(sv_x_matrix))( 7 downto 4);
                                FRM_o_B     <= E4(to_integer(sv_y_matrix),to_integer(sv_x_matrix))( 3 downto 0);
                            end if;
                            --FRM_o_R <= E4(to_integer(sv_y_matrix),to_integer(sv_x_matrix))(11 downto 8);
                            --FRM_o_G <= E4(to_integer(sv_y_matrix),to_integer(sv_x_matrix))( 7 downto 4);
                            --FRM_o_B <= E4(to_integer(sv_y_matrix),to_integer(sv_x_matrix))( 3 downto 0);
                        end if;
                        --E5
                        if ((sv_v_cnt >= 240 and sv_v_cnt <= 259 and sv_h_cnt >= 380 and sv_h_cnt <= 439) 
                            or (sv_v_cnt >= 260 and sv_v_cnt <= 279 and sv_h_cnt >= 380 and sv_h_cnt <= 399) 
                            or (sv_v_cnt >= 260 and sv_v_cnt <= 279 and sv_h_cnt >= 420 and sv_h_cnt <= 439) 
                            or (sv_v_cnt >= 280 and sv_v_cnt <= 299 and sv_h_cnt >= 380 and sv_h_cnt <= 439)) then
                            FRM_o_R <= "0000";
                            FRM_o_G <= "0000";
                            FRM_o_B <= "0000";
                        elsif (sv_v_cnt >= 260 and sv_v_cnt <= 279 and sv_h_cnt >= 400 and sv_h_cnt <= 419) then
                            sv_x_matrix <= sv_h_cnt - 400;
                            sv_y_matrix <= sv_v_cnt - 260;
                            if (si_curs_x = 5 and si_curs_y = 4) then
                                st_lamp_off <= E5;
                                FRM_o_R     <= st_cursore(to_integer(sv_y_matrix),to_integer(sv_x_matrix))(11 downto 8);
                                FRM_o_G     <= st_cursore(to_integer(sv_y_matrix),to_integer(sv_x_matrix))( 7 downto 4);
                                FRM_o_B     <= st_cursore(to_integer(sv_y_matrix),to_integer(sv_x_matrix))( 3 downto 0);
                            else
                                FRM_o_R     <= E5(to_integer(sv_y_matrix),to_integer(sv_x_matrix))(11 downto 8);
                                FRM_o_G     <= E5(to_integer(sv_y_matrix),to_integer(sv_x_matrix))( 7 downto 4);
                                FRM_o_B     <= E5(to_integer(sv_y_matrix),to_integer(sv_x_matrix))( 3 downto 0);
                            end if;
                            --FRM_o_R <= E5(to_integer(sv_y_matrix),to_integer(sv_x_matrix))(11 downto 8);
                            --FRM_o_G <= E5(to_integer(sv_y_matrix),to_integer(sv_x_matrix))( 7 downto 4);
                            --FRM_o_B <= E5(to_integer(sv_y_matrix),to_integer(sv_x_matrix))( 3 downto 0);
                        end if;
                        --E6
                        if ((sv_v_cnt >= 240 and sv_v_cnt <= 259 and sv_h_cnt >= 440 and sv_h_cnt <= 499) 
                            or (sv_v_cnt >= 260 and sv_v_cnt <= 279 and sv_h_cnt >= 440 and sv_h_cnt <= 459) 
                            or (sv_v_cnt >= 260 and sv_v_cnt <= 279 and sv_h_cnt >= 480 and sv_h_cnt <= 499) 
                            or (sv_v_cnt >= 280 and sv_v_cnt <= 299 and sv_h_cnt >= 440 and sv_h_cnt <= 499)) then
                            FRM_o_R <= "1111";
                            FRM_o_G <= "1111";
                            FRM_o_B <= "1111";
                        elsif (sv_v_cnt >= 260 and sv_v_cnt <= 279 and sv_h_cnt >= 460 and sv_h_cnt <= 479) then
                            sv_x_matrix <= sv_h_cnt - 460;
                            sv_y_matrix <= sv_v_cnt - 260;
                            if (si_curs_x = 6 and si_curs_y = 4) then
                                st_lamp_off <= E6;
                                FRM_o_R     <= st_cursore(to_integer(sv_y_matrix),to_integer(sv_x_matrix))(11 downto 8);
                                FRM_o_G     <= st_cursore(to_integer(sv_y_matrix),to_integer(sv_x_matrix))( 7 downto 4);
                                FRM_o_B     <= st_cursore(to_integer(sv_y_matrix),to_integer(sv_x_matrix))( 3 downto 0);
                            else
                                FRM_o_R     <= E6(to_integer(sv_y_matrix),to_integer(sv_x_matrix))(11 downto 8);
                                FRM_o_G     <= E6(to_integer(sv_y_matrix),to_integer(sv_x_matrix))( 7 downto 4);
                                FRM_o_B     <= E6(to_integer(sv_y_matrix),to_integer(sv_x_matrix))( 3 downto 0);
                            end if;
                            --FRM_o_R <= E6(to_integer(sv_y_matrix),to_integer(sv_x_matrix))(11 downto 8);
                            --FRM_o_G <= E6(to_integer(sv_y_matrix),to_integer(sv_x_matrix))( 7 downto 4);
                            --FRM_o_B <= E6(to_integer(sv_y_matrix),to_integer(sv_x_matrix))( 3 downto 0);
                        end if;
                        --E7
                        if ((sv_v_cnt >= 240 and sv_v_cnt <= 259 and sv_h_cnt >= 500 and sv_h_cnt <= 559) 
                            or (sv_v_cnt >= 260 and sv_v_cnt <= 279 and sv_h_cnt >= 500 and sv_h_cnt <= 519) 
                            or (sv_v_cnt >= 260 and sv_v_cnt <= 279 and sv_h_cnt >= 540 and sv_h_cnt <= 559) 
                            or (sv_v_cnt >= 280 and sv_v_cnt <= 299 and sv_h_cnt >= 500 and sv_h_cnt <= 559)) then
                            FRM_o_R <= "0000";
                            FRM_o_G <= "0000";
                            FRM_o_B <= "0000";
                        elsif (sv_v_cnt >= 260 and sv_v_cnt <= 279 and sv_h_cnt >= 520 and sv_h_cnt <= 539) then
                            sv_x_matrix <= sv_h_cnt - 520;
                            sv_y_matrix <= sv_v_cnt - 260;
                            if (si_curs_x = 7 and si_curs_y = 4) then
                                st_lamp_off <= E7;
                                FRM_o_R     <= st_cursore(to_integer(sv_y_matrix),to_integer(sv_x_matrix))(11 downto 8);
                                FRM_o_G     <= st_cursore(to_integer(sv_y_matrix),to_integer(sv_x_matrix))( 7 downto 4);
                                FRM_o_B     <= st_cursore(to_integer(sv_y_matrix),to_integer(sv_x_matrix))( 3 downto 0);
                            else
                                FRM_o_R     <= E7(to_integer(sv_y_matrix),to_integer(sv_x_matrix))(11 downto 8);
                                FRM_o_G     <= E7(to_integer(sv_y_matrix),to_integer(sv_x_matrix))( 7 downto 4);
                                FRM_o_B     <= E7(to_integer(sv_y_matrix),to_integer(sv_x_matrix))( 3 downto 0);
                            end if;
                            --FRM_o_R <= E7(to_integer(sv_y_matrix),to_integer(sv_x_matrix))(11 downto 8);
                            --FRM_o_G <= E7(to_integer(sv_y_matrix),to_integer(sv_x_matrix))( 7 downto 4);
                            --FRM_o_B <= E7(to_integer(sv_y_matrix),to_integer(sv_x_matrix))( 3 downto 0);
                        end if;
                        --F0
                        if ((sv_v_cnt >= 300 and sv_v_cnt <= 319 and sv_h_cnt >= 80 and sv_h_cnt <= 139) 
                            or (sv_v_cnt >= 320 and sv_v_cnt <= 339 and sv_h_cnt >= 80 and sv_h_cnt <= 99) 
                            or (sv_v_cnt >= 320 and sv_v_cnt <= 339 and sv_h_cnt >= 120 and sv_h_cnt <= 139) 
                            or (sv_v_cnt >= 340 and sv_v_cnt <= 359 and sv_h_cnt >= 80 and sv_h_cnt <= 139)) then
                            FRM_o_R <= "0000";
                            FRM_o_G <= "0000";
                            FRM_o_B <= "0000";
                        elsif (sv_v_cnt >= 320 and sv_v_cnt <= 339 and sv_h_cnt >= 100 and sv_h_cnt <= 119) then
                            sv_x_matrix <= sv_h_cnt - 100;
                            sv_y_matrix <= sv_v_cnt - 320;
                            if (si_curs_x = 0 and si_curs_y = 5) then
                                st_lamp_off <= F0;
                                FRM_o_R     <= st_cursore(to_integer(sv_y_matrix),to_integer(sv_x_matrix))(11 downto 8);
                                FRM_o_G     <= st_cursore(to_integer(sv_y_matrix),to_integer(sv_x_matrix))( 7 downto 4);
                                FRM_o_B     <= st_cursore(to_integer(sv_y_matrix),to_integer(sv_x_matrix))( 3 downto 0);
                            else
                                FRM_o_R     <= F0(to_integer(sv_y_matrix),to_integer(sv_x_matrix))(11 downto 8);
                                FRM_o_G     <= F0(to_integer(sv_y_matrix),to_integer(sv_x_matrix))( 7 downto 4);
                                FRM_o_B     <= F0(to_integer(sv_y_matrix),to_integer(sv_x_matrix))( 3 downto 0);
                            end if;
                            --FRM_o_R <= F0(to_integer(sv_y_matrix),to_integer(sv_x_matrix))(11 downto 8);
                            --FRM_o_G <= F0(to_integer(sv_y_matrix),to_integer(sv_x_matrix))( 7 downto 4);
                            --FRM_o_B <= F0(to_integer(sv_y_matrix),to_integer(sv_x_matrix))( 3 downto 0);
                        end if;
                        --F1
                        if ((sv_v_cnt >= 300 and sv_v_cnt <= 319 and sv_h_cnt >= 140 and sv_h_cnt <= 199) 
                            or (sv_v_cnt >= 320 and sv_v_cnt <= 339 and sv_h_cnt >= 140 and sv_h_cnt <= 159) 
                            or (sv_v_cnt >= 320 and sv_v_cnt <= 339 and sv_h_cnt >= 180 and sv_h_cnt <= 199) 
                            or (sv_v_cnt >= 340 and sv_v_cnt <= 359 and sv_h_cnt >= 140 and sv_h_cnt <= 199)) then
                            FRM_o_R <= "1111";
                            FRM_o_G <= "1111";
                            FRM_o_B <= "1111";
                        elsif (sv_v_cnt >= 320 and sv_v_cnt <= 339 and sv_h_cnt >= 160 and sv_h_cnt <= 179) then
                            sv_x_matrix <= sv_h_cnt - 160;
                            sv_y_matrix <= sv_v_cnt - 320;
                            if (si_curs_x = 1 and si_curs_y = 5) then
                                st_lamp_off <= F1;
                                FRM_o_R     <= st_cursore(to_integer(sv_y_matrix),to_integer(sv_x_matrix))(11 downto 8);
                                FRM_o_G     <= st_cursore(to_integer(sv_y_matrix),to_integer(sv_x_matrix))( 7 downto 4);
                                FRM_o_B     <= st_cursore(to_integer(sv_y_matrix),to_integer(sv_x_matrix))( 3 downto 0);
                            else
                                FRM_o_R     <= F1(to_integer(sv_y_matrix),to_integer(sv_x_matrix))(11 downto 8);
                                FRM_o_G     <= F1(to_integer(sv_y_matrix),to_integer(sv_x_matrix))( 7 downto 4);
                                FRM_o_B     <= F1(to_integer(sv_y_matrix),to_integer(sv_x_matrix))( 3 downto 0);
                            end if;
                            --FRM_o_R <= F1(to_integer(sv_y_matrix),to_integer(sv_x_matrix))(11 downto 8);
                            --FRM_o_G <= F1(to_integer(sv_y_matrix),to_integer(sv_x_matrix))( 7 downto 4);
                            --FRM_o_B <= F1(to_integer(sv_y_matrix),to_integer(sv_x_matrix))( 3 downto 0);
                        end if;
                        --F2
                        if ((sv_v_cnt >= 300 and sv_v_cnt <= 319 and sv_h_cnt >= 200 and sv_h_cnt <= 259) 
                            or (sv_v_cnt >= 320 and sv_v_cnt <= 339 and sv_h_cnt >= 200 and sv_h_cnt <= 219) 
                            or (sv_v_cnt >= 320 and sv_v_cnt <= 339 and sv_h_cnt >= 240 and sv_h_cnt <= 259) 
                            or (sv_v_cnt >= 340 and sv_v_cnt <= 359 and sv_h_cnt >= 200 and sv_h_cnt <= 259)) then
                            FRM_o_R <= "0000";
                            FRM_o_G <= "0000";
                            FRM_o_B <= "0000";
                        elsif (sv_v_cnt >= 320 and sv_v_cnt <= 339 and sv_h_cnt >= 220 and sv_h_cnt <= 239) then
                            sv_x_matrix <= sv_h_cnt - 220;
                            sv_y_matrix <= sv_v_cnt - 320;
                            if (si_curs_x = 2 and si_curs_y = 5) then
                                st_lamp_off <= F2;
                                FRM_o_R     <= st_cursore(to_integer(sv_y_matrix),to_integer(sv_x_matrix))(11 downto 8);
                                FRM_o_G     <= st_cursore(to_integer(sv_y_matrix),to_integer(sv_x_matrix))( 7 downto 4);
                                FRM_o_B     <= st_cursore(to_integer(sv_y_matrix),to_integer(sv_x_matrix))( 3 downto 0);
                            else
                                FRM_o_R     <= F2(to_integer(sv_y_matrix),to_integer(sv_x_matrix))(11 downto 8);
                                FRM_o_G     <= F2(to_integer(sv_y_matrix),to_integer(sv_x_matrix))( 7 downto 4);
                                FRM_o_B     <= F2(to_integer(sv_y_matrix),to_integer(sv_x_matrix))( 3 downto 0);
                            end if;
                            --FRM_o_R <= F2(to_integer(sv_y_matrix),to_integer(sv_x_matrix))(11 downto 8);
                            --FRM_o_G <= F2(to_integer(sv_y_matrix),to_integer(sv_x_matrix))( 7 downto 4);
                            --FRM_o_B <= F2(to_integer(sv_y_matrix),to_integer(sv_x_matrix))( 3 downto 0);
                        end if;
                        --F3
                        if ((sv_v_cnt >= 300 and sv_v_cnt <= 319 and sv_h_cnt >= 260 and sv_h_cnt <= 319) 
                            or (sv_v_cnt >= 320 and sv_v_cnt <= 339 and sv_h_cnt >= 260 and sv_h_cnt <= 279) 
                            or (sv_v_cnt >= 320 and sv_v_cnt <= 339 and sv_h_cnt >= 300 and sv_h_cnt <= 319) 
                            or (sv_v_cnt >= 340 and sv_v_cnt <= 359 and sv_h_cnt >= 260 and sv_h_cnt <= 319)) then
                            FRM_o_R <= "1111";
                            FRM_o_G <= "1111";
                            FRM_o_B <= "1111";
                        elsif (sv_v_cnt >= 320 and sv_v_cnt <= 339 and sv_h_cnt >= 280 and sv_h_cnt <= 299) then
                            sv_x_matrix <= sv_h_cnt - 280;
                            sv_y_matrix <= sv_v_cnt - 320;
                            if (si_curs_x = 3 and si_curs_y = 5) then
                                st_lamp_off <= F3;
                                FRM_o_R     <= st_cursore(to_integer(sv_y_matrix),to_integer(sv_x_matrix))(11 downto 8);
                                FRM_o_G     <= st_cursore(to_integer(sv_y_matrix),to_integer(sv_x_matrix))( 7 downto 4);
                                FRM_o_B     <= st_cursore(to_integer(sv_y_matrix),to_integer(sv_x_matrix))( 3 downto 0);
                            else
                                FRM_o_R     <= F3(to_integer(sv_y_matrix),to_integer(sv_x_matrix))(11 downto 8);
                                FRM_o_G     <= F3(to_integer(sv_y_matrix),to_integer(sv_x_matrix))( 7 downto 4);
                                FRM_o_B     <= F3(to_integer(sv_y_matrix),to_integer(sv_x_matrix))( 3 downto 0);
                            end if;
                            --FRM_o_R <= F3(to_integer(sv_y_matrix),to_integer(sv_x_matrix))(11 downto 8);
                            --FRM_o_G <= F3(to_integer(sv_y_matrix),to_integer(sv_x_matrix))( 7 downto 4);
                            --FRM_o_B <= F3(to_integer(sv_y_matrix),to_integer(sv_x_matrix))( 3 downto 0);
                        end if;
                        --F4
                        if ((sv_v_cnt >= 300 and sv_v_cnt <= 319 and sv_h_cnt >= 320 and sv_h_cnt <= 379) 
                            or (sv_v_cnt >= 320 and sv_v_cnt <= 339 and sv_h_cnt >= 320 and sv_h_cnt <= 339) 
                            or (sv_v_cnt >= 320 and sv_v_cnt <= 339 and sv_h_cnt >= 360 and sv_h_cnt <= 379) 
                            or (sv_v_cnt >= 340 and sv_v_cnt <= 359 and sv_h_cnt >= 320 and sv_h_cnt <= 379)) then
                            FRM_o_R <= "0000";
                            FRM_o_G <= "0000";
                            FRM_o_B <= "0000";
                        elsif (sv_v_cnt >= 320 and sv_v_cnt <= 339 and sv_h_cnt >= 340 and sv_h_cnt <= 359) then
                            sv_x_matrix <= sv_h_cnt - 340;
                            sv_y_matrix <= sv_v_cnt - 320;
                            if (si_curs_x = 4 and si_curs_y = 5) then
                                st_lamp_off <= F4;
                                FRM_o_R     <= st_cursore(to_integer(sv_y_matrix),to_integer(sv_x_matrix))(11 downto 8);
                                FRM_o_G     <= st_cursore(to_integer(sv_y_matrix),to_integer(sv_x_matrix))( 7 downto 4);
                                FRM_o_B     <= st_cursore(to_integer(sv_y_matrix),to_integer(sv_x_matrix))( 3 downto 0);
                            else
                                FRM_o_R     <= F4(to_integer(sv_y_matrix),to_integer(sv_x_matrix))(11 downto 8);
                                FRM_o_G     <= F4(to_integer(sv_y_matrix),to_integer(sv_x_matrix))( 7 downto 4);
                                FRM_o_B     <= F4(to_integer(sv_y_matrix),to_integer(sv_x_matrix))( 3 downto 0);
                            end if;
                            --FRM_o_R <= F4(to_integer(sv_y_matrix),to_integer(sv_x_matrix))(11 downto 8);
                            --FRM_o_G <= F4(to_integer(sv_y_matrix),to_integer(sv_x_matrix))( 7 downto 4);
                            --FRM_o_B <= F4(to_integer(sv_y_matrix),to_integer(sv_x_matrix))( 3 downto 0);
                        end if;
                        --F5
                        if ((sv_v_cnt >= 300 and sv_v_cnt <= 319 and sv_h_cnt >= 380 and sv_h_cnt <= 439) 
                            or (sv_v_cnt >= 320 and sv_v_cnt <= 339 and sv_h_cnt >= 380 and sv_h_cnt <= 399) 
                            or (sv_v_cnt >= 320 and sv_v_cnt <= 339 and sv_h_cnt >= 420 and sv_h_cnt <= 439) 
                            or (sv_v_cnt >= 340 and sv_v_cnt <= 359 and sv_h_cnt >= 380 and sv_h_cnt <= 439)) then
                            FRM_o_R <= "1111";
                            FRM_o_G <= "1111";
                            FRM_o_B <= "1111";
                        elsif (sv_v_cnt >= 320 and sv_v_cnt <= 339 and sv_h_cnt >= 400 and sv_h_cnt <= 419) then
                            sv_x_matrix <= sv_h_cnt - 400;
                            sv_y_matrix <= sv_v_cnt - 320;
                            if (si_curs_x = 5 and si_curs_y = 5) then
                                st_lamp_off <= F5;
                                FRM_o_R     <= st_cursore(to_integer(sv_y_matrix),to_integer(sv_x_matrix))(11 downto 8);
                                FRM_o_G     <= st_cursore(to_integer(sv_y_matrix),to_integer(sv_x_matrix))( 7 downto 4);
                                FRM_o_B     <= st_cursore(to_integer(sv_y_matrix),to_integer(sv_x_matrix))( 3 downto 0);
                            else
                                FRM_o_R     <= F5(to_integer(sv_y_matrix),to_integer(sv_x_matrix))(11 downto 8);
                                FRM_o_G     <= F5(to_integer(sv_y_matrix),to_integer(sv_x_matrix))( 7 downto 4);
                                FRM_o_B     <= F5(to_integer(sv_y_matrix),to_integer(sv_x_matrix))( 3 downto 0);
                            end if;
                            --FRM_o_R <= F5(to_integer(sv_y_matrix),to_integer(sv_x_matrix))(11 downto 8);
                            --FRM_o_G <= F5(to_integer(sv_x_matrix),to_integer(sv_x_matrix))( 7 downto 4);
                            --FRM_o_B <= F5(to_integer(sv_y_matrix),to_integer(sv_x_matrix))( 3 downto 0);
                        end if;
                        --F6
                        if ((sv_v_cnt >= 300 and sv_v_cnt <= 319 and sv_h_cnt >= 440 and sv_h_cnt <= 499) 
                            or (sv_v_cnt >= 320 and sv_v_cnt <= 339 and sv_h_cnt >= 440 and sv_h_cnt <= 459) 
                            or (sv_v_cnt >= 320 and sv_v_cnt <= 339 and sv_h_cnt >= 480 and sv_h_cnt <= 499) 
                            or (sv_v_cnt >= 340 and sv_v_cnt <= 359 and sv_h_cnt >= 440 and sv_h_cnt <= 499)) then
                            FRM_o_R <= "0000";
                            FRM_o_G <= "0000";
                            FRM_o_B <= "0000";
                        elsif (sv_v_cnt >= 320 and sv_v_cnt <= 339 and sv_h_cnt >= 460 and sv_h_cnt <= 479) then
                            sv_x_matrix <= sv_h_cnt - 460;
                            sv_y_matrix <= sv_v_cnt - 320;
                            if (si_curs_x = 6 and si_curs_y = 5) then
                                st_lamp_off <= F6;
                                FRM_o_R     <= st_cursore(to_integer(sv_y_matrix),to_integer(sv_x_matrix))(11 downto 8);
                                FRM_o_G     <= st_cursore(to_integer(sv_y_matrix),to_integer(sv_x_matrix))( 7 downto 4);
                                FRM_o_B     <= st_cursore(to_integer(sv_y_matrix),to_integer(sv_x_matrix))( 3 downto 0);
                            else
                                FRM_o_R     <= F6(to_integer(sv_y_matrix),to_integer(sv_x_matrix))(11 downto 8);
                                FRM_o_G     <= F6(to_integer(sv_y_matrix),to_integer(sv_x_matrix))( 7 downto 4);
                                FRM_o_B     <= F6(to_integer(sv_y_matrix),to_integer(sv_x_matrix))( 3 downto 0);
                            end if;
                            --FRM_o_R <= F6(to_integer(sv_y_matrix),to_integer(sv_x_matrix))(11 downto 8);
                            --FRM_o_G <= F6(to_integer(sv_y_matrix),to_integer(sv_x_matrix))( 7 downto 4);
                            --FRM_o_B <= F6(to_integer(sv_y_matrix),to_integer(sv_x_matrix))( 3 downto 0);
                        end if;
                        --F7
                        if ((sv_v_cnt >= 300 and sv_v_cnt <= 319 and sv_h_cnt >= 500 and sv_h_cnt <= 559) 
                            or (sv_v_cnt >= 320 and sv_v_cnt <= 339 and sv_h_cnt >= 500 and sv_h_cnt <= 519) 
                            or (sv_v_cnt >= 320 and sv_v_cnt <= 339 and sv_h_cnt >= 540 and sv_h_cnt <= 559) 
                            or (sv_v_cnt >= 340 and sv_v_cnt <= 359 and sv_h_cnt >= 500 and sv_h_cnt <= 559)) then
                            FRM_o_R <= "1111";
                            FRM_o_G <= "1111";
                            FRM_o_B <= "1111";
                        elsif (sv_v_cnt >= 320 and sv_v_cnt <= 339 and sv_h_cnt >= 520 and sv_h_cnt <= 539) then
                            sv_x_matrix <= sv_h_cnt - 520;
                            sv_y_matrix <= sv_v_cnt - 320;
                            if (si_curs_x = 7 and si_curs_y = 5) then
                                st_lamp_off <= F7;
                                FRM_o_R     <= st_cursore(to_integer(sv_y_matrix),to_integer(sv_x_matrix))(11 downto 8);
                                FRM_o_G     <= st_cursore(to_integer(sv_y_matrix),to_integer(sv_x_matrix))( 7 downto 4);
                                FRM_o_B     <= st_cursore(to_integer(sv_y_matrix),to_integer(sv_x_matrix))( 3 downto 0);
                            else
                                FRM_o_R     <= F7(to_integer(sv_y_matrix),to_integer(sv_x_matrix))(11 downto 8);
                                FRM_o_G     <= F7(to_integer(sv_y_matrix),to_integer(sv_x_matrix))( 7 downto 4);
                                FRM_o_B     <= F7(to_integer(sv_y_matrix),to_integer(sv_x_matrix))( 3 downto 0);
                            end if;
                            --FRM_o_R <= F7(to_integer(sv_y_matrix),to_integer(sv_x_matrix))(11 downto 8);
                            --FRM_o_G <= F7(to_integer(sv_y_matrix),to_integer(sv_x_matrix))( 7 downto 4);
                            --FRM_o_B <= F7(to_integer(sv_y_matrix),to_integer(sv_x_matrix))( 3 downto 0);
                        end if;
                        --G0
                        if ((sv_v_cnt >= 360 and sv_v_cnt <= 379 and sv_h_cnt >= 80 and sv_h_cnt <= 139) 
                            or (sv_v_cnt >= 380 and sv_v_cnt <= 399 and sv_h_cnt >= 80 and sv_h_cnt <= 99) 
                            or (sv_v_cnt >= 380 and sv_v_cnt <= 399 and sv_h_cnt >= 120 and sv_h_cnt <= 139) 
                            or (sv_v_cnt >= 400 and sv_v_cnt <= 419 and sv_h_cnt >= 80 and sv_h_cnt <= 139)) then
                            FRM_o_R <= "1111";
                            FRM_o_G <= "1111";
                            FRM_o_B <= "1111";
                        elsif (sv_v_cnt >= 380 and sv_v_cnt <= 399 and sv_h_cnt >= 100 and sv_h_cnt <= 119) then
                            sv_x_matrix <= sv_h_cnt - 100;
                            sv_y_matrix <= sv_v_cnt - 380;
                            if (si_curs_x = 0 and si_curs_y = 6) then
                                st_lamp_off <= G0;
                                FRM_o_R     <= st_cursore(to_integer(sv_y_matrix),to_integer(sv_x_matrix))(11 downto 8);
                                FRM_o_G     <= st_cursore(to_integer(sv_y_matrix),to_integer(sv_x_matrix))( 7 downto 4);
                                FRM_o_B     <= st_cursore(to_integer(sv_y_matrix),to_integer(sv_x_matrix))( 3 downto 0);
                            else
                                FRM_o_R     <= G0(to_integer(sv_y_matrix),to_integer(sv_x_matrix))(11 downto 8);
                                FRM_o_G     <= G0(to_integer(sv_y_matrix),to_integer(sv_x_matrix))( 7 downto 4);
                                FRM_o_B     <= G0(to_integer(sv_y_matrix),to_integer(sv_x_matrix))( 3 downto 0);
                            end if;
                            --FRM_o_R <= G0(to_integer(sv_y_matrix),to_integer(sv_x_matrix))(11 downto 8);
                            --FRM_o_G <= G0(to_integer(sv_y_matrix),to_integer(sv_x_matrix))( 7 downto 4);
                            --FRM_o_B <= G0(to_integer(sv_y_matrix),to_integer(sv_x_matrix))( 3 downto 0);
                        end if;
                        --G1
                        if ((sv_v_cnt >= 360 and sv_v_cnt <= 379 and sv_h_cnt >= 140 and sv_h_cnt <= 199) 
                            or (sv_v_cnt >= 380 and sv_v_cnt <= 399 and sv_h_cnt >= 140 and sv_h_cnt <= 159) 
                            or (sv_v_cnt >= 380 and sv_v_cnt <= 399 and sv_h_cnt >= 180 and sv_h_cnt <= 199) 
                            or (sv_v_cnt >= 400 and sv_v_cnt <= 419 and sv_h_cnt >= 140 and sv_h_cnt <= 199)) then
                            FRM_o_R <= "0000";
                            FRM_o_G <= "0000";
                            FRM_o_B <= "0000";
                        elsif (sv_v_cnt >= 380 and sv_v_cnt <= 399 and sv_h_cnt >= 160 and sv_h_cnt <= 179) then
                            sv_x_matrix <= sv_h_cnt - 160;
                            sv_y_matrix <= sv_v_cnt - 380;
                            if (si_curs_x = 1 and si_curs_y = 6) then
                                st_lamp_off <= G1;
                                FRM_o_R     <= st_cursore(to_integer(sv_y_matrix),to_integer(sv_x_matrix))(11 downto 8);
                                FRM_o_G     <= st_cursore(to_integer(sv_y_matrix),to_integer(sv_x_matrix))( 7 downto 4);
                                FRM_o_B     <= st_cursore(to_integer(sv_y_matrix),to_integer(sv_x_matrix))( 3 downto 0);
                            else
                                FRM_o_R     <= G1(to_integer(sv_y_matrix),to_integer(sv_x_matrix))(11 downto 8);
                                FRM_o_G     <= G1(to_integer(sv_y_matrix),to_integer(sv_x_matrix))( 7 downto 4);
                                FRM_o_B     <= G1(to_integer(sv_y_matrix),to_integer(sv_x_matrix))( 3 downto 0);
                            end if;
                            --FRM_o_R <= G1(to_integer(sv_y_matrix),to_integer(sv_x_matrix))(11 downto 8);
                            --FRM_o_G <= G1(to_integer(sv_y_matrix),to_integer(sv_x_matrix))( 7 downto 4);
                            --FRM_o_B <= G1(to_integer(sv_y_matrix),to_integer(sv_x_matrix))( 3 downto 0);
                        end if;
                        --G2
                        if ((sv_v_cnt >= 360 and sv_v_cnt <= 379 and sv_h_cnt >= 200 and sv_h_cnt <= 259) 
                            or (sv_v_cnt >= 380 and sv_v_cnt <= 399 and sv_h_cnt >= 200 and sv_h_cnt <= 219) 
                            or (sv_v_cnt >= 380 and sv_v_cnt <= 399 and sv_h_cnt >= 240 and sv_h_cnt <= 259) 
                            or (sv_v_cnt >= 400 and sv_v_cnt <= 419 and sv_h_cnt >= 200 and sv_h_cnt <= 259)) then
                            FRM_o_R <= "1111";
                            FRM_o_G <= "1111";
                            FRM_o_B <= "1111";
                        elsif (sv_v_cnt >= 380 and sv_v_cnt <= 399 and sv_h_cnt >= 220 and sv_h_cnt <= 239) then
                            sv_x_matrix <= sv_h_cnt - 220;
                            sv_y_matrix <= sv_v_cnt - 380;
                            if (si_curs_x = 2 and si_curs_y = 6) then
                                st_lamp_off <= G2;
                                FRM_o_R     <= st_cursore(to_integer(sv_y_matrix),to_integer(sv_x_matrix))(11 downto 8);
                                FRM_o_G     <= st_cursore(to_integer(sv_y_matrix),to_integer(sv_x_matrix))( 7 downto 4);
                                FRM_o_B     <= st_cursore(to_integer(sv_y_matrix),to_integer(sv_x_matrix))( 3 downto 0);
                            else
                                FRM_o_R     <= G2(to_integer(sv_y_matrix),to_integer(sv_x_matrix))(11 downto 8);
                                FRM_o_G     <= G2(to_integer(sv_y_matrix),to_integer(sv_x_matrix))( 7 downto 4);
                                FRM_o_B     <= G2(to_integer(sv_y_matrix),to_integer(sv_x_matrix))( 3 downto 0);
                            end if;
                            --FRM_o_R <= G2(to_integer(sv_y_matrix),to_integer(sv_x_matrix))(11 downto 8);
                            --FRM_o_G <= G2(to_integer(sv_y_matrix),to_integer(sv_x_matrix))( 7 downto 4);
                            --FRM_o_B <= G2(to_integer(sv_y_matrix),to_integer(sv_x_matrix))( 3 downto 0);
                        end if;
                        --G3
                        if ((sv_v_cnt >= 360 and sv_v_cnt <= 379 and sv_h_cnt >= 260 and sv_h_cnt <= 319) 
                            or (sv_v_cnt >= 380 and sv_v_cnt <= 399 and sv_h_cnt >= 260 and sv_h_cnt <= 279) 
                            or (sv_v_cnt >= 380 and sv_v_cnt <= 399 and sv_h_cnt >= 300 and sv_h_cnt <= 319) 
                            or (sv_v_cnt >= 400 and sv_v_cnt <= 419 and sv_h_cnt >= 260 and sv_h_cnt <= 319)) then
                            FRM_o_R <= "0000";
                            FRM_o_G <= "0000";
                            FRM_o_B <= "0000";
                        elsif (sv_v_cnt >= 380 and sv_v_cnt <= 399 and sv_h_cnt >= 280 and sv_h_cnt <= 299) then
                            sv_x_matrix <= sv_h_cnt - 280;
                            sv_y_matrix <= sv_v_cnt - 380;
                            if (si_curs_x = 3 and si_curs_y = 6) then
                                st_lamp_off <= G3;
                                FRM_o_R     <= st_cursore(to_integer(sv_y_matrix),to_integer(sv_x_matrix))(11 downto 8);
                                FRM_o_G     <= st_cursore(to_integer(sv_y_matrix),to_integer(sv_x_matrix))( 7 downto 4);
                                FRM_o_B     <= st_cursore(to_integer(sv_y_matrix),to_integer(sv_x_matrix))( 3 downto 0);
                            else
                                FRM_o_R     <= G3(to_integer(sv_y_matrix),to_integer(sv_x_matrix))(11 downto 8);
                                FRM_o_G     <= G3(to_integer(sv_y_matrix),to_integer(sv_x_matrix))( 7 downto 4);
                                FRM_o_B     <= G3(to_integer(sv_y_matrix),to_integer(sv_x_matrix))( 3 downto 0);
                            end if;
                            --FRM_o_R <= G3(to_integer(sv_y_matrix),to_integer(sv_x_matrix))(11 downto 8);
                            --FRM_o_G <= G3(to_integer(sv_y_matrix),to_integer(sv_x_matrix))( 7 downto 4);
                            --FRM_o_B <= G3(to_integer(sv_y_matrix),to_integer(sv_x_matrix))( 3 downto 0);
                        end if;
                        --G4
                        if ((sv_v_cnt >= 360 and sv_v_cnt <= 379 and sv_h_cnt >= 320 and sv_h_cnt <= 379) 
                            or (sv_v_cnt >= 380 and sv_v_cnt <= 399 and sv_h_cnt >= 320 and sv_h_cnt <= 339) 
                            or (sv_v_cnt >= 380 and sv_v_cnt <= 399 and sv_h_cnt >= 360 and sv_h_cnt <= 379) 
                            or (sv_v_cnt >= 400 and sv_v_cnt <= 419 and sv_h_cnt >= 320 and sv_h_cnt <= 379)) then
                            FRM_o_R <= "1111";
                            FRM_o_G <= "1111";
                            FRM_o_B <= "1111";
                        elsif (sv_v_cnt >= 380 and sv_v_cnt <= 399 and sv_h_cnt >= 340 and sv_h_cnt <= 359) then
                            sv_x_matrix <= sv_h_cnt - 340;
                            sv_y_matrix <= sv_v_cnt - 380;
                            if (si_curs_x = 4 and si_curs_y = 6) then
                                st_lamp_off <= G4;
                                FRM_o_R     <= st_cursore(to_integer(sv_y_matrix),to_integer(sv_x_matrix))(11 downto 8);
                                FRM_o_G     <= st_cursore(to_integer(sv_y_matrix),to_integer(sv_x_matrix))( 7 downto 4);
                                FRM_o_B     <= st_cursore(to_integer(sv_y_matrix),to_integer(sv_x_matrix))( 3 downto 0);
                            else
                                FRM_o_R     <= G4(to_integer(sv_y_matrix),to_integer(sv_x_matrix))(11 downto 8);
                                FRM_o_G     <= G4(to_integer(sv_y_matrix),to_integer(sv_x_matrix))( 7 downto 4);
                                FRM_o_B     <= G4(to_integer(sv_y_matrix),to_integer(sv_x_matrix))( 3 downto 0);
                            end if;
                            --FRM_o_R <= G4(to_integer(sv_y_matrix),to_integer(sv_x_matrix))(11 downto 8);
                            --FRM_o_G <= G4(to_integer(sv_y_matrix),to_integer(sv_x_matrix))( 7 downto 4);
                            --FRM_o_B <= G4(to_integer(sv_y_matrix),to_integer(sv_x_matrix))( 3 downto 0);
                        end if;
                        --G5
                        if ((sv_v_cnt >= 360 and sv_v_cnt <= 379 and sv_h_cnt >= 380 and sv_h_cnt <= 439) 
                            or (sv_v_cnt >= 380 and sv_v_cnt <= 399 and sv_h_cnt >= 380 and sv_h_cnt <= 399) 
                            or (sv_v_cnt >= 380 and sv_v_cnt <= 399 and sv_h_cnt >= 420 and sv_h_cnt <= 439) 
                            or (sv_v_cnt >= 400 and sv_v_cnt <= 419 and sv_h_cnt >= 380 and sv_h_cnt <= 439)) then
                            FRM_o_R <= "0000";
                            FRM_o_G <= "0000";
                            FRM_o_B <= "0000";
                        elsif (sv_v_cnt >= 380 and sv_v_cnt <= 399 and sv_h_cnt >= 400 and sv_h_cnt <= 419) then
                            sv_x_matrix <= sv_h_cnt - 400;
                            sv_y_matrix <= sv_v_cnt - 380;
                            if (si_curs_x = 5 and si_curs_y = 6) then
                                st_lamp_off <= G5;
                                FRM_o_R     <= st_cursore(to_integer(sv_y_matrix),to_integer(sv_x_matrix))(11 downto 8);
                                FRM_o_G     <= st_cursore(to_integer(sv_y_matrix),to_integer(sv_x_matrix))( 7 downto 4);
                                FRM_o_B     <= st_cursore(to_integer(sv_y_matrix),to_integer(sv_x_matrix))( 3 downto 0);
                            else
                                FRM_o_R     <= G5(to_integer(sv_y_matrix),to_integer(sv_x_matrix))(11 downto 8);
                                FRM_o_G     <= G5(to_integer(sv_y_matrix),to_integer(sv_x_matrix))( 7 downto 4);
                                FRM_o_B     <= G5(to_integer(sv_y_matrix),to_integer(sv_x_matrix))( 3 downto 0);
                            end if;
                            --FRM_o_R <= G5(to_integer(sv_y_matrix),to_integer(sv_x_matrix))(11 downto 8);
                            --FRM_o_G <= G5(to_integer(sv_y_matrix),to_integer(sv_x_matrix))( 7 downto 4);
                            --FRM_o_B <= G5(to_integer(sv_y_matrix),to_integer(sv_x_matrix))( 3 downto 0);
                        end if;
                        --G6
                        if ((sv_v_cnt >= 360 and sv_v_cnt <= 379 and sv_h_cnt >= 440 and sv_h_cnt <= 499) 
                            or (sv_v_cnt >= 380 and sv_v_cnt <= 399 and sv_h_cnt >= 440 and sv_h_cnt <= 459) 
                            or (sv_v_cnt >= 380 and sv_v_cnt <= 399 and sv_h_cnt >= 480 and sv_h_cnt <= 499) 
                            or (sv_v_cnt >= 400 and sv_v_cnt <= 419 and sv_h_cnt >= 440 and sv_h_cnt <= 499)) then
                            FRM_o_R <= "1111";
                            FRM_o_G <= "1111";
                            FRM_o_B <= "1111";
                        elsif (sv_v_cnt >= 380 and sv_v_cnt <= 399 and sv_h_cnt >= 460 and sv_h_cnt <= 479) then
                            sv_x_matrix <= sv_h_cnt - 460;
                            sv_y_matrix <= sv_v_cnt - 380;
                            if (si_curs_x = 6 and si_curs_y = 6) then
                                st_lamp_off <= G6;
                                FRM_o_R     <= st_cursore(to_integer(sv_y_matrix),to_integer(sv_x_matrix))(11 downto 8);
                                FRM_o_G     <= st_cursore(to_integer(sv_y_matrix),to_integer(sv_x_matrix))( 7 downto 4);
                                FRM_o_B     <= st_cursore(to_integer(sv_y_matrix),to_integer(sv_x_matrix))( 3 downto 0);
                            else
                                FRM_o_R     <= G6(to_integer(sv_y_matrix),to_integer(sv_x_matrix))(11 downto 8);
                                FRM_o_G     <= G6(to_integer(sv_y_matrix),to_integer(sv_x_matrix))( 7 downto 4);
                                FRM_o_B     <= G6(to_integer(sv_y_matrix),to_integer(sv_x_matrix))( 3 downto 0);
                            end if;
                            --FRM_o_R <= G6(to_integer(sv_y_matrix),to_integer(sv_x_matrix))(11 downto 8);
                            --FRM_o_G <= G6(to_integer(sv_y_matrix),to_integer(sv_x_matrix))( 7 downto 4);
                            --FRM_o_B <= G6(to_integer(sv_y_matrix),to_integer(sv_x_matrix))( 3 downto 0);
                        end if;
                        --G7
                        if ((sv_v_cnt >= 360 and sv_v_cnt <= 379 and sv_h_cnt >= 500 and sv_h_cnt <= 559) 
                            or (sv_v_cnt >= 380 and sv_v_cnt <= 399 and sv_h_cnt >= 500 and sv_h_cnt <= 519) 
                            or (sv_v_cnt >= 380 and sv_v_cnt <= 399 and sv_h_cnt >= 540 and sv_h_cnt <= 559) 
                            or (sv_v_cnt >= 400 and sv_v_cnt <= 419 and sv_h_cnt >= 500 and sv_h_cnt <= 559)) then
                            FRM_o_R <= "0000";
                            FRM_o_G <= "0000";
                            FRM_o_B <= "0000";
                        elsif (sv_v_cnt >= 380 and sv_v_cnt <= 399 and sv_h_cnt >= 520 and sv_h_cnt <= 539) then
                            sv_x_matrix <= sv_h_cnt - 520;
                            sv_y_matrix <= sv_v_cnt - 380;
                            if (si_curs_x = 7 and si_curs_y = 6) then
                                st_lamp_off <= G7;
                                FRM_o_R     <= st_cursore(to_integer(sv_y_matrix),to_integer(sv_x_matrix))(11 downto 8);
                                FRM_o_G     <= st_cursore(to_integer(sv_y_matrix),to_integer(sv_x_matrix))( 7 downto 4);
                                FRM_o_B     <= st_cursore(to_integer(sv_y_matrix),to_integer(sv_x_matrix))( 3 downto 0);
                            else
                                FRM_o_R     <= G7(to_integer(sv_y_matrix),to_integer(sv_x_matrix))(11 downto 8);
                                FRM_o_G     <= G7(to_integer(sv_y_matrix),to_integer(sv_x_matrix))( 7 downto 4);
                                FRM_o_B     <= G7(to_integer(sv_y_matrix),to_integer(sv_x_matrix))( 3 downto 0);
                            end if;
                            --FRM_o_R <= G7(to_integer(sv_y_matrix),to_integer(sv_x_matrix))(11 downto 8);
                            --FRM_o_G <= G7(to_integer(sv_y_matrix),to_integer(sv_x_matrix))( 7 downto 4);
                            --FRM_o_B <= G7(to_integer(sv_y_matrix),to_integer(sv_x_matrix))( 3 downto 0);
                        end if;
                        --H0
                        if ((sv_v_cnt >= 420 and sv_v_cnt <= 439 and sv_h_cnt >= 80 and sv_h_cnt <= 139) 
                            or (sv_v_cnt >= 440 and sv_v_cnt <= 459 and sv_h_cnt >= 80 and sv_h_cnt <= 99) 
                            or (sv_v_cnt >= 440 and sv_v_cnt <= 459 and sv_h_cnt >= 120 and sv_h_cnt <= 139) 
                            or (sv_v_cnt >= 460 and sv_v_cnt <= 479 and sv_h_cnt >= 80 and sv_h_cnt <= 139)) then
                            FRM_o_R <= "0000";
                            FRM_o_G <= "0000";
                            FRM_o_B <= "0000";
                        elsif (sv_v_cnt >= 440 and sv_v_cnt <= 459 and sv_h_cnt >= 100 and sv_h_cnt <= 119) then
                            sv_x_matrix <= sv_h_cnt - 100;
                            sv_y_matrix <= sv_v_cnt - 440;
                            if (si_curs_x = 0 and si_curs_y = 7) then
                                st_lamp_off <= H0;
                                FRM_o_R     <= st_cursore(to_integer(sv_y_matrix),to_integer(sv_x_matrix))(11 downto 8);
                                FRM_o_G     <= st_cursore(to_integer(sv_y_matrix),to_integer(sv_x_matrix))( 7 downto 4);
                                FRM_o_B     <= st_cursore(to_integer(sv_y_matrix),to_integer(sv_x_matrix))( 3 downto 0);
                            else
                                FRM_o_R     <= H0(to_integer(sv_y_matrix),to_integer(sv_x_matrix))(11 downto 8);
                                FRM_o_G     <= H0(to_integer(sv_y_matrix),to_integer(sv_x_matrix))( 7 downto 4);
                                FRM_o_B     <= H0(to_integer(sv_y_matrix),to_integer(sv_x_matrix))( 3 downto 0);
                            end if;
                            --FRM_o_R <= H0(to_integer(sv_y_matrix),to_integer(sv_x_matrix))(11 downto 8);
                            --FRM_o_G <= H0(to_integer(sv_y_matrix),to_integer(sv_x_matrix))( 7 downto 4);
                            --FRM_o_B <= H0(to_integer(sv_y_matrix),to_integer(sv_x_matrix))( 3 downto 0);
                        end if;
                        --H1
                        if ((sv_v_cnt >= 420 and sv_v_cnt <= 439 and sv_h_cnt >= 140 and sv_h_cnt <= 199) 
                            or (sv_v_cnt >= 440 and sv_v_cnt <= 459 and sv_h_cnt >= 140 and sv_h_cnt <= 159) 
                            or (sv_v_cnt >= 440 and sv_v_cnt <= 459 and sv_h_cnt >= 180 and sv_h_cnt <= 199) 
                            or (sv_v_cnt >= 460 and sv_v_cnt <= 479 and sv_h_cnt >= 140 and sv_h_cnt <= 199)) then
                            FRM_o_R <= "1111";
                            FRM_o_G <= "1111";
                            FRM_o_B <= "1111";
                        elsif (sv_v_cnt >= 440 and sv_v_cnt <= 459 and sv_h_cnt >= 160 and sv_h_cnt <= 179) then
                            sv_x_matrix <= sv_h_cnt - 160;
                            sv_y_matrix <= sv_v_cnt - 440;
                            if (si_curs_x = 1 and si_curs_y = 7) then
                                st_lamp_off <= H1;
                                FRM_o_R     <= st_cursore(to_integer(sv_y_matrix),to_integer(sv_x_matrix))(11 downto 8);
                                FRM_o_G     <= st_cursore(to_integer(sv_y_matrix),to_integer(sv_x_matrix))( 7 downto 4);
                                FRM_o_B     <= st_cursore(to_integer(sv_y_matrix),to_integer(sv_x_matrix))( 3 downto 0);
                            else
                                FRM_o_R     <= H1(to_integer(sv_y_matrix),to_integer(sv_x_matrix))(11 downto 8);
                                FRM_o_G     <= H1(to_integer(sv_y_matrix),to_integer(sv_x_matrix))( 7 downto 4);
                                FRM_o_B     <= H1(to_integer(sv_y_matrix),to_integer(sv_x_matrix))( 3 downto 0);
                            end if;
                            --FRM_o_R <= H1(to_integer(sv_y_matrix),to_integer(sv_x_matrix))(11 downto 8);
                            --FRM_o_G <= H1(to_integer(sv_y_matrix),to_integer(sv_x_matrix))( 7 downto 4);
                            --FRM_o_B <= H1(to_integer(sv_y_matrix),to_integer(sv_x_matrix))( 3 downto 0);
                        end if;
                        --H2
                        if ((sv_v_cnt >= 420 and sv_v_cnt <= 439 and sv_h_cnt >= 200 and sv_h_cnt <= 259) 
                            or (sv_v_cnt >= 440 and sv_v_cnt <= 459 and sv_h_cnt >= 200 and sv_h_cnt <= 219) 
                            or (sv_v_cnt >= 440 and sv_v_cnt <= 459 and sv_h_cnt >= 240 and sv_h_cnt <= 259) 
                            or (sv_v_cnt >= 460 and sv_v_cnt <= 479 and sv_h_cnt >= 200 and sv_h_cnt <= 259)) then
                            FRM_o_R <= "0000";
                            FRM_o_G <= "0000";
                            FRM_o_B <= "0000";
                        elsif (sv_v_cnt >= 440 and sv_v_cnt <= 459 and sv_h_cnt >= 220 and sv_h_cnt <= 239) then
                            sv_x_matrix <= sv_h_cnt - 220;
                            sv_y_matrix <= sv_v_cnt - 440;
                            if (si_curs_x = 2 and si_curs_y = 7) then
                                st_lamp_off <= H2;
                                FRM_o_R     <= st_cursore(to_integer(sv_y_matrix),to_integer(sv_x_matrix))(11 downto 8);
                                FRM_o_G     <= st_cursore(to_integer(sv_y_matrix),to_integer(sv_x_matrix))( 7 downto 4);
                                FRM_o_B     <= st_cursore(to_integer(sv_y_matrix),to_integer(sv_x_matrix))( 3 downto 0);
                            else
                                FRM_o_R     <= H2(to_integer(sv_y_matrix),to_integer(sv_x_matrix))(11 downto 8);
                                FRM_o_G     <= H2(to_integer(sv_y_matrix),to_integer(sv_x_matrix))( 7 downto 4);
                                FRM_o_B     <= H2(to_integer(sv_y_matrix),to_integer(sv_x_matrix))( 3 downto 0);
                            end if;
                            --FRM_o_R <= H2(to_integer(sv_y_matrix),to_integer(sv_x_matrix))(11 downto 8);
                            --FRM_o_G <= H2(to_integer(sv_y_matrix),to_integer(sv_x_matrix))( 7 downto 4);
                            --FRM_o_B <= H2(to_integer(sv_y_matrix),to_integer(sv_x_matrix))( 3 downto 0);
                        end if;
                        --H3
                        if ((sv_v_cnt >= 420 and sv_v_cnt <= 439 and sv_h_cnt >= 260 and sv_h_cnt <= 319) 
                            or (sv_v_cnt >= 440 and sv_v_cnt <= 459 and sv_h_cnt >= 260 and sv_h_cnt <= 279) 
                            or (sv_v_cnt >= 440 and sv_v_cnt <= 459 and sv_h_cnt >= 300 and sv_h_cnt <= 319) 
                            or (sv_v_cnt >= 460 and sv_v_cnt <= 479 and sv_h_cnt >= 260 and sv_h_cnt <= 319)) then
                            FRM_o_R <= "1111";
                            FRM_o_G <= "1111";
                            FRM_o_B <= "1111";
                        elsif (sv_v_cnt >= 440 and sv_v_cnt <= 459 and sv_h_cnt >= 280 and sv_h_cnt <= 299) then
                            sv_x_matrix <= sv_h_cnt - 280;
                            sv_y_matrix <= sv_v_cnt - 440;
                            if (si_curs_x = 3 and si_curs_y = 7) then
                                st_lamp_off <= H3;
                                FRM_o_R     <= st_cursore(to_integer(sv_y_matrix),to_integer(sv_x_matrix))(11 downto 8);
                                FRM_o_G     <= st_cursore(to_integer(sv_y_matrix),to_integer(sv_x_matrix))( 7 downto 4);
                                FRM_o_B     <= st_cursore(to_integer(sv_y_matrix),to_integer(sv_x_matrix))( 3 downto 0);
                            else
                                FRM_o_R     <= H3(to_integer(sv_y_matrix),to_integer(sv_x_matrix))(11 downto 8);
                                FRM_o_G     <= H3(to_integer(sv_y_matrix),to_integer(sv_x_matrix))( 7 downto 4);
                                FRM_o_B     <= H3(to_integer(sv_y_matrix),to_integer(sv_x_matrix))( 3 downto 0);
                            end if;
                            --FRM_o_R <= H3(to_integer(sv_y_matrix),to_integer(sv_x_matrix))(11 downto 8);
                            --FRM_o_G <= H3(to_integer(sv_y_matrix),to_integer(sv_x_matrix))( 7 downto 4);
                            --FRM_o_B <= H3(to_integer(sv_y_matrix),to_integer(sv_x_matrix))( 3 downto 0);
                        end if;
                        --H4
                        if ((sv_v_cnt >= 420 and sv_v_cnt <= 439 and sv_h_cnt >= 320 and sv_h_cnt <= 379) 
                            or (sv_v_cnt >= 440 and sv_v_cnt <= 459 and sv_h_cnt >= 320 and sv_h_cnt <= 339) 
                            or (sv_v_cnt >= 440 and sv_v_cnt <= 459 and sv_h_cnt >= 360 and sv_h_cnt <= 379) 
                            or (sv_v_cnt >= 460 and sv_v_cnt <= 479 and sv_h_cnt >= 320 and sv_h_cnt <= 379)) then
                            FRM_o_R <= "0000";
                            FRM_o_G <= "0000";
                            FRM_o_B <= "0000";
                        elsif (sv_v_cnt >= 440 and sv_v_cnt <= 459 and sv_h_cnt >= 340 and sv_h_cnt <= 359) then
                            sv_x_matrix <= sv_h_cnt - 340;
                            sv_y_matrix <= sv_v_cnt - 440;
                            if (si_curs_x = 4 and si_curs_y = 7) then
                                st_lamp_off <= H4;
                                FRM_o_R     <= st_cursore(to_integer(sv_y_matrix),to_integer(sv_x_matrix))(11 downto 8);
                                FRM_o_G     <= st_cursore(to_integer(sv_y_matrix),to_integer(sv_x_matrix))( 7 downto 4);
                                FRM_o_B     <= st_cursore(to_integer(sv_y_matrix),to_integer(sv_x_matrix))( 3 downto 0);
                            else
                                FRM_o_R     <= H4(to_integer(sv_y_matrix),to_integer(sv_x_matrix))(11 downto 8);
                                FRM_o_G     <= H4(to_integer(sv_y_matrix),to_integer(sv_x_matrix))( 7 downto 4);
                                FRM_o_B     <= H4(to_integer(sv_y_matrix),to_integer(sv_x_matrix))( 3 downto 0);
                            end if;
                            --FRM_o_R <= H4(to_integer(sv_y_matrix),to_integer(sv_x_matrix))(11 downto 8);
                            --FRM_o_G <= H4(to_integer(sv_y_matrix),to_integer(sv_x_matrix))( 7 downto 4);
                            --FRM_o_B <= H4(to_integer(sv_y_matrix),to_integer(sv_x_matrix))( 3 downto 0);
                        end if;
                        --H5
                        if ((sv_v_cnt >= 420 and sv_v_cnt <= 439 and sv_h_cnt >= 380 and sv_h_cnt <= 439) 
                            or (sv_v_cnt >= 440 and sv_v_cnt <= 459 and sv_h_cnt >= 380 and sv_h_cnt <= 399) 
                            or (sv_v_cnt >= 440 and sv_v_cnt <= 459 and sv_h_cnt >= 420 and sv_h_cnt <= 439) 
                            or (sv_v_cnt >= 460 and sv_v_cnt <= 479 and sv_h_cnt >= 380 and sv_h_cnt <= 439)) then
                            FRM_o_R <= "1111";
                            FRM_o_G <= "1111";
                            FRM_o_B <= "1111";
                        elsif (sv_v_cnt >= 440 and sv_v_cnt <= 459 and sv_h_cnt >= 400 and sv_h_cnt <= 419) then
                            sv_x_matrix <= sv_h_cnt - 400;
                            sv_y_matrix <= sv_v_cnt - 440;
                            if (si_curs_x = 5 and si_curs_y = 7) then
                                st_lamp_off <= H5;
                                FRM_o_R     <= st_cursore(to_integer(sv_y_matrix),to_integer(sv_x_matrix))(11 downto 8);
                                FRM_o_G     <= st_cursore(to_integer(sv_y_matrix),to_integer(sv_x_matrix))( 7 downto 4);
                                FRM_o_B     <= st_cursore(to_integer(sv_y_matrix),to_integer(sv_x_matrix))( 3 downto 0);
                            else
                                FRM_o_R     <= H5(to_integer(sv_y_matrix),to_integer(sv_x_matrix))(11 downto 8);
                                FRM_o_G     <= H5(to_integer(sv_y_matrix),to_integer(sv_x_matrix))( 7 downto 4);
                                FRM_o_B     <= H5(to_integer(sv_y_matrix),to_integer(sv_x_matrix))( 3 downto 0);
                            end if;
                            --FRM_o_R <= H5(to_integer(sv_y_matrix),to_integer(sv_x_matrix))(11 downto 8);
                            --FRM_o_G <= H5(to_integer(sv_y_matrix),to_integer(sv_x_matrix))( 7 downto 4);
                            --FRM_o_B <= H5(to_integer(sv_y_matrix),to_integer(sv_x_matrix))( 3 downto 0);
                        end if;
                        --H6
                        if ((sv_v_cnt >= 420 and sv_v_cnt <= 439 and sv_h_cnt >= 440 and sv_h_cnt <= 499) 
                            or (sv_v_cnt >= 440 and sv_v_cnt <= 459 and sv_h_cnt >= 440 and sv_h_cnt <= 459) 
                            or (sv_v_cnt >= 440 and sv_v_cnt <= 459 and sv_h_cnt >= 480 and sv_h_cnt <= 499) 
                            or (sv_v_cnt >= 460 and sv_v_cnt <= 479 and sv_h_cnt >= 440 and sv_h_cnt <= 499)) then
                            FRM_o_R <= "0000";
                            FRM_o_G <= "0000";
                            FRM_o_B <= "0000";
                        elsif (sv_v_cnt >= 440 and sv_v_cnt <= 459 and sv_h_cnt >= 460 and sv_h_cnt <= 479) then
                            sv_x_matrix <= sv_h_cnt - 460;
                            sv_y_matrix <= sv_v_cnt - 440;
                            if (si_curs_x = 6 and si_curs_y = 7) then
                                st_lamp_off <= H6;
                                FRM_o_R     <= st_cursore(to_integer(sv_y_matrix),to_integer(sv_x_matrix))(11 downto 8);
                                FRM_o_G     <= st_cursore(to_integer(sv_y_matrix),to_integer(sv_x_matrix))( 7 downto 4);
                                FRM_o_B     <= st_cursore(to_integer(sv_y_matrix),to_integer(sv_x_matrix))( 3 downto 0);
                            else
                                FRM_o_R     <= H6(to_integer(sv_y_matrix),to_integer(sv_x_matrix))(11 downto 8);
                                FRM_o_G     <= H6(to_integer(sv_y_matrix),to_integer(sv_x_matrix))( 7 downto 4);
                                FRM_o_B     <= H6(to_integer(sv_y_matrix),to_integer(sv_x_matrix))( 3 downto 0);
                            end if;
                            --FRM_o_R <= H6(to_integer(sv_y_matrix),to_integer(sv_x_matrix))(11 downto 8);
                            --FRM_o_G <= H6(to_integer(sv_y_matrix),to_integer(sv_x_matrix))( 7 downto 4);
                            --FRM_o_B <= H6(to_integer(sv_y_matrix),to_integer(sv_x_matrix))( 3 downto 0);
                        end if;
                        --H7
                        if ((sv_v_cnt >= 420 and sv_v_cnt <= 439 and sv_h_cnt >= 500 and sv_h_cnt <= 559) 
                            or (sv_v_cnt >= 440 and sv_v_cnt <= 459 and sv_h_cnt >= 500 and sv_h_cnt <= 519) 
                            or (sv_v_cnt >= 440 and sv_v_cnt <= 459 and sv_h_cnt >= 540 and sv_h_cnt <= 559) 
                            or (sv_v_cnt >= 460 and sv_v_cnt <= 479 and sv_h_cnt >= 500 and sv_h_cnt <= 559)) then
                            FRM_o_R <= "1111";
                            FRM_o_G <= "1111";
                            FRM_o_B <= "1111";
                        elsif (sv_v_cnt >= 440 and sv_v_cnt <= 459 and sv_h_cnt >= 520 and sv_h_cnt <= 539) then
                            sv_x_matrix <= sv_h_cnt - 520;
                            sv_y_matrix <= sv_v_cnt - 440;
                            if (si_curs_x = 7 and si_curs_y = 7) then
                                st_lamp_off <= H7;
                                FRM_o_R     <= st_cursore(to_integer(sv_y_matrix),to_integer(sv_x_matrix))(11 downto 8);
                                FRM_o_G     <= st_cursore(to_integer(sv_y_matrix),to_integer(sv_x_matrix))( 7 downto 4);
                                FRM_o_B     <= st_cursore(to_integer(sv_y_matrix),to_integer(sv_x_matrix))( 3 downto 0);
                            else
                                FRM_o_R     <= H7(to_integer(sv_y_matrix),to_integer(sv_x_matrix))(11 downto 8);
                                FRM_o_G     <= H7(to_integer(sv_y_matrix),to_integer(sv_x_matrix))( 7 downto 4);
                                FRM_o_B     <= H7(to_integer(sv_y_matrix),to_integer(sv_x_matrix))( 3 downto 0);
                            end if;
                            --FRM_o_R <= H7(to_integer(sv_y_matrix),to_integer(sv_x_matrix))(11 downto 8);
                            --FRM_o_G <= H7(to_integer(sv_y_matrix),to_integer(sv_x_matrix))( 7 downto 4);
                            --FRM_o_B <= H7(to_integer(sv_y_matrix),to_integer(sv_x_matrix))( 3 downto 0);
                        end if;
                        --fuori
                        if ((sv_h_cnt >= 0 and sv_h_cnt <= 79) or (sv_h_cnt >= 560 and sv_h_cnt <= 639)) then --grigio scuro: 010001000100
                            FRM_o_R <= "0100";  
                            FRM_o_G <= "0100";
                            FRM_o_B <= "0100";
                        end if;            
                    end if;
            end if;
        end process;
                     
end Behavioral;
